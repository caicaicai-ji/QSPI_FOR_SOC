/*
     Copyright (c) 2018 SMIC             
     Filename:      qspi_info_fifo_mem.lef
     IP code:       S55NLLG2PH
     Version:       1.1.0
     CreateDate:    Oct 31, 2018        
                    
    LEF for General 2-PORT SRAM
    SMIC 55nm LL Logic Process

    Configuration: -instname qspi_info_fifo_mem -rows 32 -bits 16 -mux 1 
    Redundancy: Off
    Bit-Write: Off
*/

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO qspi_info_fifo_mem
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 100.74 BY 58.915 ;

 PIN QA[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[0]

 PIN QA[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[1]

 PIN QA[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[2]

 PIN QA[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[3]

 PIN QA[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[4]

 PIN QA[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[5]

 PIN QA[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[6]

 PIN QA[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[7]

 PIN AA[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 37.055 58.915 37.255 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 37.055 58.915 37.255 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 37.055 58.915 37.255 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[1]

 PIN AA[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 40.16 58.915 40.36 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 40.16 58.915 40.36 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 40.16 58.915 40.36 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[0]

 PIN AA[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 40.81 58.915 41.01 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 40.81 58.915 41.01 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 40.81 58.915 41.01 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[2]

 PIN AA[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 46.71 58.915 46.91 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 46.71 58.915 46.91 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 46.71 58.915 46.91 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[4]

 PIN AA[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 48.145 58.915 48.345 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 48.145 58.915 48.345 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 48.145 58.915 48.345 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[3]

 PIN CENA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 73.47 58.915 73.67 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 73.47 58.915 73.67 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 73.47 58.915 73.67 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENA

 PIN CLKA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 73.96 58.915 74.16 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 73.96 58.915 74.16 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 73.96 58.915 74.16 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKA

 PIN QA[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 81.775 58.915 81.975 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 81.775 58.915 81.975 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 81.775 58.915 81.975 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[8]

 PIN QA[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 82.865 58.915 83.065 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 82.865 58.915 83.065 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 82.865 58.915 83.065 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[9]

 PIN QA[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 86.315 58.915 86.515 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 86.315 58.915 86.515 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 86.315 58.915 86.515 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[10]

 PIN QA[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 87.405 58.915 87.605 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 87.405 58.915 87.605 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 87.405 58.915 87.605 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[11]

 PIN QA[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 90.855 58.915 91.055 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 90.855 58.915 91.055 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 90.855 58.915 91.055 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[12]

 PIN QA[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 91.945 58.915 92.145 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 91.945 58.915 92.145 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 91.945 58.915 92.145 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[13]

 PIN QA[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 95.395 58.915 95.595 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 95.395 58.915 95.595 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 95.395 58.915 95.595 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[14]

 PIN QA[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 96.485 58.915 96.685 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 96.485 58.915 96.685 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 96.485 58.915 96.685 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[15]

 PIN DB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[0]

 PIN DB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[1]

 PIN DB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[2]

 PIN DB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[3]

 PIN DB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[4]

 PIN DB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[5]

 PIN DB[6]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[6]

 PIN DB[7]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[7]

 PIN CLKB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.85 0 24.05 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.85 0 24.05 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.85 0 24.05 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKB

 PIN CENB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 24.34 0 24.54 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 24.34 0 24.54 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 24.34 0 24.54 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENB

 PIN AB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 49.44 0 49.64 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 49.44 0 49.64 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 49.44 0 49.64 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[3]

 PIN AB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 50.875 0 51.075 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 50.875 0 51.075 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 50.875 0 51.075 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[4]

 PIN AB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 56.775 0 56.975 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 56.775 0 56.975 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 56.775 0 56.975 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[2]

 PIN AB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 57.425 0 57.625 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 57.425 0 57.625 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 57.425 0 57.625 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[0]

 PIN AB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 60.53 0 60.73 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 60.53 0 60.73 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 60.53 0 60.73 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[1]

 PIN DB[8]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 81.53 0 81.73 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 81.53 0 81.73 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 81.53 0 81.73 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[8]

 PIN DB[9]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 83.11 0 83.31 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 83.11 0 83.31 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 83.11 0 83.31 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[9]

 PIN DB[10]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 86.07 0 86.27 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 86.07 0 86.27 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 86.07 0 86.27 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[10]

 PIN DB[11]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 87.65 0 87.85 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 87.65 0 87.85 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 87.65 0 87.85 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[11]

 PIN DB[12]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 90.61 0 90.81 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 90.61 0 90.81 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 90.61 0 90.81 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[12]

 PIN DB[13]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 92.19 0 92.39 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 92.19 0 92.39 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 92.19 0 92.39 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[13]

 PIN DB[14]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 95.15 0 95.35 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 95.15 0 95.35 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 95.15 0 95.35 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[14]

 PIN DB[15]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 96.73 0 96.93 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 96.73 0 96.93 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 96.73 0 96.93 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[15]

 PIN VDD
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 2.43 0 3.93 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.01 0 11.51 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 11.51 0 13.01 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 19.09 0 20.59 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 23.81 0 28.81 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 34.26 0 37.76 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 41.96 0 45.96 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 54.78 0 58.78 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 62.98 0 66.48 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 71.93 0 76.93 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 80.15 0 81.65 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 87.73 0 89.23 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 89.23 0 90.73 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 96.81 0 98.31 58.915 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 5.47 0 6.97 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 6.97 0 8.47 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 14.55 0 16.05 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 16.05 0 17.55 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 29.66 0 33.66 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 38.36 0 41.36 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 47.365 0 53.365 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 59.38 0 62.38 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 67.08 0 71.08 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 83.19 0 84.69 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 84.69 0 86.19 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 92.27 0 93.77 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 93.77 0 95.27 58.915 ;      
 END
 END VSS

 OBS
 LAYER M1 ;
 RECT 0 0 3.72 0.585 ;
 RECT 4.1 0 5.3 0.585 ;
 RECT 5.68 0 8.26 0.585 ;
 RECT 8.64 0 9.84 0.585 ;
 RECT 10.22 0 12.8 0.585 ;
 RECT 13.18 0 14.38 0.585 ;
 RECT 14.76 0 17.34 0.585 ;
 RECT 17.72 0 18.92 0.585 ;
 RECT 19.3 0 23.76 0.585 ;
 RECT 24.14 0 24.25 0.585 ;
 RECT 24.63 0 49.35 0.585 ;
 RECT 49.73 0 50.785 0.585 ;
 RECT 51.165 0 56.685 0.585 ;
 RECT 57.065 0 57.335 0.585 ;
 RECT 57.715 0 60.44 0.585 ;
 RECT 60.82 0 81.44 0.585 ;
 RECT 81.82 0 83.02 0.585 ;
 RECT 83.4 0 85.98 0.585 ;
 RECT 86.36 0 87.56 0.585 ;
 RECT 87.94 0 90.52 0.585 ;
 RECT 90.9 0 92.1 0.585 ;
 RECT 92.48 0 95.06 0.585 ;
 RECT 95.44 0 96.64 0.585 ;
 RECT 97.02 0 100.74 0.585 ;
 RECT 0 58.915 3.965 58.33 ;
 RECT 4.345 58.915 5.055 58.33 ;
 RECT 5.435 58.915 8.505 58.33 ;
 RECT 8.885 58.915 9.595 58.33 ;
 RECT 9.975 58.915 13.045 58.33 ;
 RECT 13.425 58.915 14.135 58.33 ;
 RECT 14.515 58.915 17.585 58.33 ;
 RECT 17.965 58.915 18.675 58.33 ;
 RECT 19.055 58.915 36.965 58.33 ;
 RECT 37.345 58.915 40.07 58.33 ;
 RECT 40.45 58.915 40.72 58.33 ;
 RECT 41.1 58.915 46.62 58.33 ;
 RECT 47 58.915 48.055 58.33 ;
 RECT 48.435 58.915 73.38 58.33 ;
 RECT 73.76 58.915 73.87 58.33 ;
 RECT 74.25 58.915 81.685 58.33 ;
 RECT 82.065 58.915 82.775 58.33 ;
 RECT 83.155 58.915 86.225 58.33 ;
 RECT 86.605 58.915 87.315 58.33 ;
 RECT 87.695 58.915 90.765 58.33 ;
 RECT 91.145 58.915 91.855 58.33 ;
 RECT 92.235 58.915 95.305 58.33 ;
 RECT 95.685 58.915 96.395 58.33 ;
 RECT 96.775 58.915 100.74 58.33 ;
 RECT 0 0.585 100.74 58.33 ;
 LAYER M2 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 23.75 0.595 ;
 RECT 24.64 0 49.34 0.595 ;
 RECT 49.74 0 50.775 0.595 ;
 RECT 51.175 0 56.675 0.595 ;
 RECT 57.075 0 57.325 0.595 ;
 RECT 57.725 0 60.43 0.595 ;
 RECT 60.83 0 81.43 0.595 ;
 RECT 81.83 0 83.01 0.595 ;
 RECT 83.41 0 85.97 0.595 ;
 RECT 86.37 0 87.55 0.595 ;
 RECT 87.95 0 90.51 0.595 ;
 RECT 90.91 0 92.09 0.595 ;
 RECT 92.49 0 95.05 0.595 ;
 RECT 95.45 0 96.63 0.595 ;
 RECT 97.03 0 100.74 0.595 ;
 RECT 0 58.915 3.955 58.32 ;
 RECT 4.355 58.915 5.045 58.32 ;
 RECT 5.445 58.915 8.495 58.32 ;
 RECT 8.895 58.915 9.585 58.32 ;
 RECT 9.985 58.915 13.035 58.32 ;
 RECT 13.435 58.915 14.125 58.32 ;
 RECT 14.525 58.915 17.575 58.32 ;
 RECT 17.975 58.915 18.665 58.32 ;
 RECT 19.065 58.915 36.955 58.32 ;
 RECT 37.355 58.915 40.06 58.32 ;
 RECT 40.46 58.915 40.71 58.32 ;
 RECT 41.11 58.915 46.61 58.32 ;
 RECT 47.01 58.915 48.045 58.32 ;
 RECT 48.445 58.915 73.37 58.32 ;
 RECT 74.26 58.915 81.675 58.32 ;
 RECT 82.075 58.915 82.765 58.32 ;
 RECT 83.165 58.915 86.215 58.32 ;
 RECT 86.615 58.915 87.305 58.32 ;
 RECT 87.705 58.915 90.755 58.32 ;
 RECT 91.155 58.915 91.845 58.32 ;
 RECT 92.245 58.915 95.295 58.32 ;
 RECT 95.695 58.915 96.385 58.32 ;
 RECT 96.785 58.915 100.74 58.32 ;
 RECT 0 0.595 100.74 58.32 ;
 LAYER M3 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 23.75 0.595 ;
 RECT 24.64 0 49.34 0.595 ;
 RECT 49.74 0 50.775 0.595 ;
 RECT 51.175 0 56.675 0.595 ;
 RECT 57.075 0 57.325 0.595 ;
 RECT 57.725 0 60.43 0.595 ;
 RECT 60.83 0 81.43 0.595 ;
 RECT 81.83 0 83.01 0.595 ;
 RECT 83.41 0 85.97 0.595 ;
 RECT 86.37 0 87.55 0.595 ;
 RECT 87.95 0 90.51 0.595 ;
 RECT 90.91 0 92.09 0.595 ;
 RECT 92.49 0 95.05 0.595 ;
 RECT 95.45 0 96.63 0.595 ;
 RECT 97.03 0 100.74 0.595 ;
 RECT 0 58.915 3.955 58.32 ;
 RECT 4.355 58.915 5.045 58.32 ;
 RECT 5.445 58.915 8.495 58.32 ;
 RECT 8.895 58.915 9.585 58.32 ;
 RECT 9.985 58.915 13.035 58.32 ;
 RECT 13.435 58.915 14.125 58.32 ;
 RECT 14.525 58.915 17.575 58.32 ;
 RECT 17.975 58.915 18.665 58.32 ;
 RECT 19.065 58.915 36.955 58.32 ;
 RECT 37.355 58.915 40.06 58.32 ;
 RECT 40.46 58.915 40.71 58.32 ;
 RECT 41.11 58.915 46.61 58.32 ;
 RECT 47.01 58.915 48.045 58.32 ;
 RECT 48.445 58.915 73.37 58.32 ;
 RECT 74.26 58.915 81.675 58.32 ;
 RECT 82.075 58.915 82.765 58.32 ;
 RECT 83.165 58.915 86.215 58.32 ;
 RECT 86.615 58.915 87.305 58.32 ;
 RECT 87.705 58.915 90.755 58.32 ;
 RECT 91.155 58.915 91.845 58.32 ;
 RECT 92.245 58.915 95.295 58.32 ;
 RECT 95.695 58.915 96.385 58.32 ;
 RECT 96.785 58.915 100.74 58.32 ;
 RECT 0 0.595 100.74 58.32 ;

 LAYER V1 ;
 RECT 0 0 100.74 58.915 ;
 LAYER V2 ;
 RECT 0 0 100.74 58.915 ;
 LAYER V3 ;
 RECT 0 0 100.74 58.915 ;

 LAYER M4 ;
 RECT 20.69 0 23.71 0.595 ;
 RECT 20.69 0.595 23.71 58.915 ;
 RECT 28.91 0 29.56 0.595 ;
 RECT 28.91 0.595 29.56 58.915 ;
 RECT 33.76 0 34.16 0.595 ;
 RECT 33.76 0.595 34.16 58.915 ;
 RECT 37.86 0 38.26 0.595 ;
 RECT 37.86 0.595 38.26 58.915 ;
 RECT 41.46 0 41.86 0.595 ;
 RECT 41.46 0.595 41.86 58.915 ;
 RECT 46.06 0 47.265 0.595 ;
 RECT 46.06 0.595 47.265 58.915 ;
 RECT 53.465 0 54.68 0.595 ;
 RECT 53.465 0.595 54.68 58.915 ;
 RECT 58.88 0 59.28 0.595 ;
 RECT 58.88 0.595 59.28 58.915 ;
 RECT 62.48 0 62.88 0.595 ;
 RECT 62.48 0.595 62.88 58.915 ;
 RECT 66.58 0 66.98 0.595 ;
 RECT 66.58 0.595 66.98 58.915 ;
 RECT 71.18 0 71.83 0.595 ;
 RECT 71.18 0.595 71.83 58.915 ;
 RECT 77.03 0 80.05 0.595 ;
 RECT 77.03 0.595 80.05 58.915 ;
 LAYER V4 ;
 RECT 20.69 0 23.71 0.595 ;
 RECT 20.69 0.595 23.71 58.915 ;
 RECT 28.91 0 29.56 0.595 ;
 RECT 28.91 0.595 29.56 58.915 ;
 RECT 33.76 0 34.16 0.595 ;
 RECT 33.76 0.595 34.16 58.915 ;
 RECT 37.86 0 38.26 0.595 ;
 RECT 37.86 0.595 38.26 58.915 ;
 RECT 41.46 0 41.86 0.595 ;
 RECT 41.46 0.595 41.86 58.915 ;
 RECT 46.06 0 47.265 0.595 ;
 RECT 46.06 0.595 47.265 58.915 ;
 RECT 53.465 0 54.68 0.595 ;
 RECT 53.465 0.595 54.68 58.915 ;
 RECT 58.88 0 59.28 0.595 ;
 RECT 58.88 0.595 59.28 58.915 ;
 RECT 62.48 0 62.88 0.595 ;
 RECT 62.48 0.595 62.88 58.915 ;
 RECT 66.58 0 66.98 0.595 ;
 RECT 66.58 0.595 66.98 58.915 ;
 RECT 71.18 0 71.83 0.595 ;
 RECT 71.18 0.595 71.83 58.915 ;
 RECT 77.03 0 80.05 0.595 ;
 RECT 77.03 0.595 80.05 58.915 ;
 END

END qspi_info_fifo_mem
END LIBRARY