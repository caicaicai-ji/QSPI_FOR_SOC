/*
     Copyright (c) 2018 SMIC             
     Filename:      qspi_addr_fifo_mem.lef
     IP code:       S55NLLG2PH
     Version:       1.1.0
     CreateDate:    Oct 31, 2018        
                    
    LEF for General 2-PORT SRAM
    SMIC 55nm LL Logic Process

    Configuration: -instname qspi_addr_fifo_mem -rows 32 -bits 32 -mux 1 
    Redundancy: Off
    Bit-Write: Off
*/

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO qspi_addr_fifo_mem
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 137.06 BY 58.915 ;

 PIN QA[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 4.055 58.915 4.255 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[0]

 PIN QA[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.145 58.915 5.345 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[1]

 PIN QA[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.595 58.915 8.795 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[2]

 PIN QA[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.685 58.915 9.885 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[3]

 PIN QA[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 13.135 58.915 13.335 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[4]

 PIN QA[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.225 58.915 14.425 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[5]

 PIN QA[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.675 58.915 17.875 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[6]

 PIN QA[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 18.765 58.915 18.965 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[7]

 PIN QA[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 22.215 58.915 22.415 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 22.215 58.915 22.415 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 22.215 58.915 22.415 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[8]

 PIN QA[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.305 58.915 23.505 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.305 58.915 23.505 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.305 58.915 23.505 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[9]

 PIN QA[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.755 58.915 26.955 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.755 58.915 26.955 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.755 58.915 26.955 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[10]

 PIN QA[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 27.845 58.915 28.045 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 27.845 58.915 28.045 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 27.845 58.915 28.045 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[11]

 PIN QA[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.295 58.915 31.495 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.295 58.915 31.495 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.295 58.915 31.495 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[12]

 PIN QA[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.385 58.915 32.585 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.385 58.915 32.585 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.385 58.915 32.585 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[13]

 PIN QA[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.835 58.915 36.035 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.835 58.915 36.035 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.835 58.915 36.035 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[14]

 PIN QA[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 36.925 58.915 37.125 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 36.925 58.915 37.125 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 36.925 58.915 37.125 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[15]

 PIN AA[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 55.215 58.915 55.415 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 55.215 58.915 55.415 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 55.215 58.915 55.415 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[1]

 PIN AA[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.32 58.915 58.52 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.32 58.915 58.52 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.32 58.915 58.52 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[0]

 PIN AA[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.97 58.915 59.17 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.97 58.915 59.17 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.97 58.915 59.17 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[2]

 PIN AA[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 64.87 58.915 65.07 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 64.87 58.915 65.07 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 64.87 58.915 65.07 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[4]

 PIN AA[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 66.305 58.915 66.505 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 66.305 58.915 66.505 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 66.305 58.915 66.505 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[3]

 PIN CENA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 91.63 58.915 91.83 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 91.63 58.915 91.83 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 91.63 58.915 91.83 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENA

 PIN CLKA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 92.12 58.915 92.32 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 92.12 58.915 92.32 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 92.12 58.915 92.32 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKA

 PIN QA[16]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 99.935 58.915 100.135 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 99.935 58.915 100.135 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 99.935 58.915 100.135 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[16]

 PIN QA[17]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 101.025 58.915 101.225 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 101.025 58.915 101.225 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 101.025 58.915 101.225 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[17]

 PIN QA[18]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 104.475 58.915 104.675 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 104.475 58.915 104.675 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 104.475 58.915 104.675 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[18]

 PIN QA[19]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 105.565 58.915 105.765 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 105.565 58.915 105.765 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 105.565 58.915 105.765 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[19]

 PIN QA[20]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 109.015 58.915 109.215 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 109.015 58.915 109.215 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 109.015 58.915 109.215 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[20]

 PIN QA[21]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 110.105 58.915 110.305 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 110.105 58.915 110.305 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 110.105 58.915 110.305 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[21]

 PIN QA[22]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 113.555 58.915 113.755 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 113.555 58.915 113.755 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 113.555 58.915 113.755 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[22]

 PIN QA[23]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 114.645 58.915 114.845 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 114.645 58.915 114.845 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 114.645 58.915 114.845 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[23]

 PIN QA[24]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 118.095 58.915 118.295 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 118.095 58.915 118.295 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 118.095 58.915 118.295 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[24]

 PIN QA[25]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 119.185 58.915 119.385 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 119.185 58.915 119.385 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 119.185 58.915 119.385 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[25]

 PIN QA[26]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 122.635 58.915 122.835 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 122.635 58.915 122.835 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 122.635 58.915 122.835 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[26]

 PIN QA[27]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 123.725 58.915 123.925 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 123.725 58.915 123.925 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 123.725 58.915 123.925 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[27]

 PIN QA[28]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 127.175 58.915 127.375 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 127.175 58.915 127.375 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 127.175 58.915 127.375 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[28]

 PIN QA[29]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 128.265 58.915 128.465 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 128.265 58.915 128.465 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 128.265 58.915 128.465 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[29]

 PIN QA[30]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 131.715 58.915 131.915 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 131.715 58.915 131.915 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 131.715 58.915 131.915 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[30]

 PIN QA[31]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 132.805 58.915 133.005 58.42 ;
 END
 PORT
 LAYER M2 ;
 RECT 132.805 58.915 133.005 58.42 ;
 END
 PORT
 LAYER M1 ;
 RECT 132.805 58.915 133.005 58.42 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[31]

 PIN DB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[0]

 PIN DB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[1]

 PIN DB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[2]

 PIN DB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[3]

 PIN DB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[4]

 PIN DB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[5]

 PIN DB[6]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[6]

 PIN DB[7]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[7]

 PIN DB[8]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[8]

 PIN DB[9]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[9]

 PIN DB[10]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[10]

 PIN DB[11]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[11]

 PIN DB[12]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[12]

 PIN DB[13]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[13]

 PIN DB[14]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[14]

 PIN DB[15]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[15]

 PIN CLKB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKB

 PIN CENB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENB

 PIN AB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[3]

 PIN AB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[4]

 PIN AB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[2]

 PIN AB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[0]

 PIN AB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[1]

 PIN DB[16]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[16]

 PIN DB[17]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[17]

 PIN DB[18]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[18]

 PIN DB[19]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[19]

 PIN DB[20]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[20]

 PIN DB[21]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[21]

 PIN DB[22]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[22]

 PIN DB[23]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[23]

 PIN DB[24]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[24]

 PIN DB[25]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[25]

 PIN DB[26]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[26]

 PIN DB[27]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[27]

 PIN DB[28]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[28]

 PIN DB[29]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[29]

 PIN DB[30]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[30]

 PIN DB[31]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[31]

 PIN VDD
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 2.43 0 3.93 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.01 0 11.51 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 11.51 0 13.01 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 19.09 0 20.59 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 20.59 0 22.09 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 28.17 0 29.67 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 29.67 0 31.17 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 37.25 0 38.75 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 41.97 0 46.97 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 52.42 0 55.92 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 60.12 0 64.12 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 72.94 0 76.94 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 81.14 0 84.64 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 90.09 0 95.09 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 98.31 0 99.81 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 105.89 0 107.39 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 107.39 0 108.89 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 114.97 0 116.47 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 116.47 0 117.97 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 124.05 0 125.55 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 125.55 0 127.05 58.915 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 133.13 0 134.63 58.915 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 5.47 0 6.97 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 6.97 0 8.47 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 14.55 0 16.05 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 16.05 0 17.55 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 23.63 0 25.13 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 25.13 0 26.63 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 32.71 0 34.21 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 34.21 0 35.71 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 47.82 0 51.82 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 56.52 0 59.52 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 65.525 0 71.525 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 77.54 0 80.54 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 85.24 0 89.24 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 101.35 0 102.85 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 102.85 0 104.35 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 110.43 0 111.93 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 111.93 0 113.43 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 119.51 0 121.01 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 121.01 0 122.51 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 128.59 0 130.09 58.915 ;      
 END
 PORT
 LAYER M4 ;
 RECT 130.09 0 131.59 58.915 ;      
 END
 END VSS

 OBS
 LAYER M1 ;
 RECT 0 0 3.72 0.585 ;
 RECT 4.1 0 5.3 0.585 ;
 RECT 5.68 0 8.26 0.585 ;
 RECT 8.64 0 9.84 0.585 ;
 RECT 10.22 0 12.8 0.585 ;
 RECT 13.18 0 14.38 0.585 ;
 RECT 14.76 0 17.34 0.585 ;
 RECT 17.72 0 18.92 0.585 ;
 RECT 19.3 0 21.88 0.585 ;
 RECT 22.26 0 23.46 0.585 ;
 RECT 23.84 0 26.42 0.585 ;
 RECT 26.8 0 28 0.585 ;
 RECT 28.38 0 30.96 0.585 ;
 RECT 31.34 0 32.54 0.585 ;
 RECT 32.92 0 35.5 0.585 ;
 RECT 35.88 0 37.08 0.585 ;
 RECT 37.46 0 41.92 0.585 ;
 RECT 42.3 0 42.41 0.585 ;
 RECT 42.79 0 67.51 0.585 ;
 RECT 67.89 0 68.945 0.585 ;
 RECT 69.325 0 74.845 0.585 ;
 RECT 75.225 0 75.495 0.585 ;
 RECT 75.875 0 78.6 0.585 ;
 RECT 78.98 0 99.6 0.585 ;
 RECT 99.98 0 101.18 0.585 ;
 RECT 101.56 0 104.14 0.585 ;
 RECT 104.52 0 105.72 0.585 ;
 RECT 106.1 0 108.68 0.585 ;
 RECT 109.06 0 110.26 0.585 ;
 RECT 110.64 0 113.22 0.585 ;
 RECT 113.6 0 114.8 0.585 ;
 RECT 115.18 0 117.76 0.585 ;
 RECT 118.14 0 119.34 0.585 ;
 RECT 119.72 0 122.3 0.585 ;
 RECT 122.68 0 123.88 0.585 ;
 RECT 124.26 0 126.84 0.585 ;
 RECT 127.22 0 128.42 0.585 ;
 RECT 128.8 0 131.38 0.585 ;
 RECT 131.76 0 132.96 0.585 ;
 RECT 133.34 0 137.06 0.585 ;
 RECT 0 58.915 3.965 58.33 ;
 RECT 4.345 58.915 5.055 58.33 ;
 RECT 5.435 58.915 8.505 58.33 ;
 RECT 8.885 58.915 9.595 58.33 ;
 RECT 9.975 58.915 13.045 58.33 ;
 RECT 13.425 58.915 14.135 58.33 ;
 RECT 14.515 58.915 17.585 58.33 ;
 RECT 17.965 58.915 18.675 58.33 ;
 RECT 19.055 58.915 22.125 58.33 ;
 RECT 22.505 58.915 23.215 58.33 ;
 RECT 23.595 58.915 26.665 58.33 ;
 RECT 27.045 58.915 27.755 58.33 ;
 RECT 28.135 58.915 31.205 58.33 ;
 RECT 31.585 58.915 32.295 58.33 ;
 RECT 32.675 58.915 35.745 58.33 ;
 RECT 36.125 58.915 36.835 58.33 ;
 RECT 37.215 58.915 55.125 58.33 ;
 RECT 55.505 58.915 58.23 58.33 ;
 RECT 58.61 58.915 58.88 58.33 ;
 RECT 59.26 58.915 64.78 58.33 ;
 RECT 65.16 58.915 66.215 58.33 ;
 RECT 66.595 58.915 91.54 58.33 ;
 RECT 91.92 58.915 92.03 58.33 ;
 RECT 92.41 58.915 99.845 58.33 ;
 RECT 100.225 58.915 100.935 58.33 ;
 RECT 101.315 58.915 104.385 58.33 ;
 RECT 104.765 58.915 105.475 58.33 ;
 RECT 105.855 58.915 108.925 58.33 ;
 RECT 109.305 58.915 110.015 58.33 ;
 RECT 110.395 58.915 113.465 58.33 ;
 RECT 113.845 58.915 114.555 58.33 ;
 RECT 114.935 58.915 118.005 58.33 ;
 RECT 118.385 58.915 119.095 58.33 ;
 RECT 119.475 58.915 122.545 58.33 ;
 RECT 122.925 58.915 123.635 58.33 ;
 RECT 124.015 58.915 127.085 58.33 ;
 RECT 127.465 58.915 128.175 58.33 ;
 RECT 128.555 58.915 131.625 58.33 ;
 RECT 132.005 58.915 132.715 58.33 ;
 RECT 133.095 58.915 137.06 58.33 ;
 RECT 0 0.585 137.06 58.33 ;
 LAYER M2 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 41.91 0.595 ;
 RECT 42.8 0 67.5 0.595 ;
 RECT 67.9 0 68.935 0.595 ;
 RECT 69.335 0 74.835 0.595 ;
 RECT 75.235 0 75.485 0.595 ;
 RECT 75.885 0 78.59 0.595 ;
 RECT 78.99 0 99.59 0.595 ;
 RECT 99.99 0 101.17 0.595 ;
 RECT 101.57 0 104.13 0.595 ;
 RECT 104.53 0 105.71 0.595 ;
 RECT 106.11 0 108.67 0.595 ;
 RECT 109.07 0 110.25 0.595 ;
 RECT 110.65 0 113.21 0.595 ;
 RECT 113.61 0 114.79 0.595 ;
 RECT 115.19 0 117.75 0.595 ;
 RECT 118.15 0 119.33 0.595 ;
 RECT 119.73 0 122.29 0.595 ;
 RECT 122.69 0 123.87 0.595 ;
 RECT 124.27 0 126.83 0.595 ;
 RECT 127.23 0 128.41 0.595 ;
 RECT 128.81 0 131.37 0.595 ;
 RECT 131.77 0 132.95 0.595 ;
 RECT 133.35 0 137.06 0.595 ;
 RECT 0 58.915 3.955 58.32 ;
 RECT 4.355 58.915 5.045 58.32 ;
 RECT 5.445 58.915 8.495 58.32 ;
 RECT 8.895 58.915 9.585 58.32 ;
 RECT 9.985 58.915 13.035 58.32 ;
 RECT 13.435 58.915 14.125 58.32 ;
 RECT 14.525 58.915 17.575 58.32 ;
 RECT 17.975 58.915 18.665 58.32 ;
 RECT 19.065 58.915 22.115 58.32 ;
 RECT 22.515 58.915 23.205 58.32 ;
 RECT 23.605 58.915 26.655 58.32 ;
 RECT 27.055 58.915 27.745 58.32 ;
 RECT 28.145 58.915 31.195 58.32 ;
 RECT 31.595 58.915 32.285 58.32 ;
 RECT 32.685 58.915 35.735 58.32 ;
 RECT 36.135 58.915 36.825 58.32 ;
 RECT 37.225 58.915 55.115 58.32 ;
 RECT 55.515 58.915 58.22 58.32 ;
 RECT 58.62 58.915 58.87 58.32 ;
 RECT 59.27 58.915 64.77 58.32 ;
 RECT 65.17 58.915 66.205 58.32 ;
 RECT 66.605 58.915 91.53 58.32 ;
 RECT 92.42 58.915 99.835 58.32 ;
 RECT 100.235 58.915 100.925 58.32 ;
 RECT 101.325 58.915 104.375 58.32 ;
 RECT 104.775 58.915 105.465 58.32 ;
 RECT 105.865 58.915 108.915 58.32 ;
 RECT 109.315 58.915 110.005 58.32 ;
 RECT 110.405 58.915 113.455 58.32 ;
 RECT 113.855 58.915 114.545 58.32 ;
 RECT 114.945 58.915 117.995 58.32 ;
 RECT 118.395 58.915 119.085 58.32 ;
 RECT 119.485 58.915 122.535 58.32 ;
 RECT 122.935 58.915 123.625 58.32 ;
 RECT 124.025 58.915 127.075 58.32 ;
 RECT 127.475 58.915 128.165 58.32 ;
 RECT 128.565 58.915 131.615 58.32 ;
 RECT 132.015 58.915 132.705 58.32 ;
 RECT 133.105 58.915 137.06 58.32 ;
 RECT 0 0.595 137.06 58.32 ;
 LAYER M3 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 41.91 0.595 ;
 RECT 42.8 0 67.5 0.595 ;
 RECT 67.9 0 68.935 0.595 ;
 RECT 69.335 0 74.835 0.595 ;
 RECT 75.235 0 75.485 0.595 ;
 RECT 75.885 0 78.59 0.595 ;
 RECT 78.99 0 99.59 0.595 ;
 RECT 99.99 0 101.17 0.595 ;
 RECT 101.57 0 104.13 0.595 ;
 RECT 104.53 0 105.71 0.595 ;
 RECT 106.11 0 108.67 0.595 ;
 RECT 109.07 0 110.25 0.595 ;
 RECT 110.65 0 113.21 0.595 ;
 RECT 113.61 0 114.79 0.595 ;
 RECT 115.19 0 117.75 0.595 ;
 RECT 118.15 0 119.33 0.595 ;
 RECT 119.73 0 122.29 0.595 ;
 RECT 122.69 0 123.87 0.595 ;
 RECT 124.27 0 126.83 0.595 ;
 RECT 127.23 0 128.41 0.595 ;
 RECT 128.81 0 131.37 0.595 ;
 RECT 131.77 0 132.95 0.595 ;
 RECT 133.35 0 137.06 0.595 ;
 RECT 0 58.915 3.955 58.32 ;
 RECT 4.355 58.915 5.045 58.32 ;
 RECT 5.445 58.915 8.495 58.32 ;
 RECT 8.895 58.915 9.585 58.32 ;
 RECT 9.985 58.915 13.035 58.32 ;
 RECT 13.435 58.915 14.125 58.32 ;
 RECT 14.525 58.915 17.575 58.32 ;
 RECT 17.975 58.915 18.665 58.32 ;
 RECT 19.065 58.915 22.115 58.32 ;
 RECT 22.515 58.915 23.205 58.32 ;
 RECT 23.605 58.915 26.655 58.32 ;
 RECT 27.055 58.915 27.745 58.32 ;
 RECT 28.145 58.915 31.195 58.32 ;
 RECT 31.595 58.915 32.285 58.32 ;
 RECT 32.685 58.915 35.735 58.32 ;
 RECT 36.135 58.915 36.825 58.32 ;
 RECT 37.225 58.915 55.115 58.32 ;
 RECT 55.515 58.915 58.22 58.32 ;
 RECT 58.62 58.915 58.87 58.32 ;
 RECT 59.27 58.915 64.77 58.32 ;
 RECT 65.17 58.915 66.205 58.32 ;
 RECT 66.605 58.915 91.53 58.32 ;
 RECT 92.42 58.915 99.835 58.32 ;
 RECT 100.235 58.915 100.925 58.32 ;
 RECT 101.325 58.915 104.375 58.32 ;
 RECT 104.775 58.915 105.465 58.32 ;
 RECT 105.865 58.915 108.915 58.32 ;
 RECT 109.315 58.915 110.005 58.32 ;
 RECT 110.405 58.915 113.455 58.32 ;
 RECT 113.855 58.915 114.545 58.32 ;
 RECT 114.945 58.915 117.995 58.32 ;
 RECT 118.395 58.915 119.085 58.32 ;
 RECT 119.485 58.915 122.535 58.32 ;
 RECT 122.935 58.915 123.625 58.32 ;
 RECT 124.025 58.915 127.075 58.32 ;
 RECT 127.475 58.915 128.165 58.32 ;
 RECT 128.565 58.915 131.615 58.32 ;
 RECT 132.015 58.915 132.705 58.32 ;
 RECT 133.105 58.915 137.06 58.32 ;
 RECT 0 0.595 137.06 58.32 ;

 LAYER V1 ;
 RECT 0 0 137.06 58.915 ;
 LAYER V2 ;
 RECT 0 0 137.06 58.915 ;
 LAYER V3 ;
 RECT 0 0 137.06 58.915 ;

 LAYER M4 ;
 RECT 38.85 0 41.87 0.595 ;
 RECT 38.85 0.595 41.87 58.915 ;
 RECT 47.07 0 47.72 0.595 ;
 RECT 47.07 0.595 47.72 58.915 ;
 RECT 51.92 0 52.32 0.595 ;
 RECT 51.92 0.595 52.32 58.915 ;
 RECT 56.02 0 56.42 0.595 ;
 RECT 56.02 0.595 56.42 58.915 ;
 RECT 59.62 0 60.02 0.595 ;
 RECT 59.62 0.595 60.02 58.915 ;
 RECT 64.22 0 65.425 0.595 ;
 RECT 64.22 0.595 65.425 58.915 ;
 RECT 71.625 0 72.84 0.595 ;
 RECT 71.625 0.595 72.84 58.915 ;
 RECT 77.04 0 77.44 0.595 ;
 RECT 77.04 0.595 77.44 58.915 ;
 RECT 80.64 0 81.04 0.595 ;
 RECT 80.64 0.595 81.04 58.915 ;
 RECT 84.74 0 85.14 0.595 ;
 RECT 84.74 0.595 85.14 58.915 ;
 RECT 89.34 0 89.99 0.595 ;
 RECT 89.34 0.595 89.99 58.915 ;
 RECT 95.19 0 98.21 0.595 ;
 RECT 95.19 0.595 98.21 58.915 ;
 LAYER V4 ;
 RECT 38.85 0 41.87 0.595 ;
 RECT 38.85 0.595 41.87 58.915 ;
 RECT 47.07 0 47.72 0.595 ;
 RECT 47.07 0.595 47.72 58.915 ;
 RECT 51.92 0 52.32 0.595 ;
 RECT 51.92 0.595 52.32 58.915 ;
 RECT 56.02 0 56.42 0.595 ;
 RECT 56.02 0.595 56.42 58.915 ;
 RECT 59.62 0 60.02 0.595 ;
 RECT 59.62 0.595 60.02 58.915 ;
 RECT 64.22 0 65.425 0.595 ;
 RECT 64.22 0.595 65.425 58.915 ;
 RECT 71.625 0 72.84 0.595 ;
 RECT 71.625 0.595 72.84 58.915 ;
 RECT 77.04 0 77.44 0.595 ;
 RECT 77.04 0.595 77.44 58.915 ;
 RECT 80.64 0 81.04 0.595 ;
 RECT 80.64 0.595 81.04 58.915 ;
 RECT 84.74 0 85.14 0.595 ;
 RECT 84.74 0.595 85.14 58.915 ;
 RECT 89.34 0 89.99 0.595 ;
 RECT 89.34 0.595 89.99 58.915 ;
 RECT 95.19 0 98.21 0.595 ;
 RECT 95.19 0.595 98.21 58.915 ;
 END

END qspi_addr_fifo_mem
END LIBRARY