/*
     Copyright (c) 2018 SMIC             
     Filename:      qspi_data_info_64_mem.lef
     IP code:       S55NLLG2PH
     Version:       1.1.0
     CreateDate:    Oct 28, 2018        
                    
    LEF for General 2-PORT SRAM
    SMIC 55nm LL Logic Process

    Configuration: -instname qspi_data_info_64_mem -rows 64 -bits 64 -mux 1 
    Redundancy: Off
    Bit-Write: Off
*/

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO qspi_data_info_64_mem
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 209.7 BY 76.575 ;

 PIN QA[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[0]

 PIN QA[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[1]

 PIN QA[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[2]

 PIN QA[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[3]

 PIN QA[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[4]

 PIN QA[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[5]

 PIN QA[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[6]

 PIN QA[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[7]

 PIN QA[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[8]

 PIN QA[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[9]

 PIN QA[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[10]

 PIN QA[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[11]

 PIN QA[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[12]

 PIN QA[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[13]

 PIN QA[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[14]

 PIN QA[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[15]

 PIN QA[16]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 40.375 76.575 40.575 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 40.375 76.575 40.575 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 40.375 76.575 40.575 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[16]

 PIN QA[17]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 41.465 76.575 41.665 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 41.465 76.575 41.665 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 41.465 76.575 41.665 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[17]

 PIN QA[18]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 44.915 76.575 45.115 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 44.915 76.575 45.115 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 44.915 76.575 45.115 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[18]

 PIN QA[19]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 46.005 76.575 46.205 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 46.005 76.575 46.205 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 46.005 76.575 46.205 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[19]

 PIN QA[20]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 49.455 76.575 49.655 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 49.455 76.575 49.655 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 49.455 76.575 49.655 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[20]

 PIN QA[21]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 50.545 76.575 50.745 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 50.545 76.575 50.745 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 50.545 76.575 50.745 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[21]

 PIN QA[22]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 53.995 76.575 54.195 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 53.995 76.575 54.195 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 53.995 76.575 54.195 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[22]

 PIN QA[23]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 55.085 76.575 55.285 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 55.085 76.575 55.285 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 55.085 76.575 55.285 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[23]

 PIN QA[24]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.535 76.575 58.735 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.535 76.575 58.735 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.535 76.575 58.735 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[24]

 PIN QA[25]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 59.625 76.575 59.825 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 59.625 76.575 59.825 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 59.625 76.575 59.825 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[25]

 PIN QA[26]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 63.075 76.575 63.275 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 63.075 76.575 63.275 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 63.075 76.575 63.275 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[26]

 PIN QA[27]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 64.165 76.575 64.365 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 64.165 76.575 64.365 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 64.165 76.575 64.365 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[27]

 PIN QA[28]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 67.615 76.575 67.815 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 67.615 76.575 67.815 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 67.615 76.575 67.815 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[28]

 PIN QA[29]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 68.705 76.575 68.905 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 68.705 76.575 68.905 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 68.705 76.575 68.905 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[29]

 PIN QA[30]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 72.155 76.575 72.355 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 72.155 76.575 72.355 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 72.155 76.575 72.355 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[30]

 PIN QA[31]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 73.245 76.575 73.445 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 73.245 76.575 73.445 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 73.245 76.575 73.445 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[31]

 PIN AA[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 91.535 76.575 91.735 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 91.535 76.575 91.735 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 91.535 76.575 91.735 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[1]

 PIN AA[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 94.64 76.575 94.84 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 94.64 76.575 94.84 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 94.64 76.575 94.84 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[0]

 PIN AA[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 95.29 76.575 95.49 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 95.29 76.575 95.49 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 95.29 76.575 95.49 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[2]

 PIN AA[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 101.19 76.575 101.39 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 101.19 76.575 101.39 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 101.19 76.575 101.39 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[4]

 PIN AA[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 102.625 76.575 102.825 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 102.625 76.575 102.825 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 102.625 76.575 102.825 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[3]

 PIN AA[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 106.115 76.575 106.315 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 106.115 76.575 106.315 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 106.115 76.575 106.315 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[5]

 PIN CENA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 127.95 76.575 128.15 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 127.95 76.575 128.15 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 127.95 76.575 128.15 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENA

 PIN CLKA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 128.44 76.575 128.64 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 128.44 76.575 128.64 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 128.44 76.575 128.64 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKA

 PIN QA[32]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 136.255 76.575 136.455 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 136.255 76.575 136.455 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 136.255 76.575 136.455 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[32]

 PIN QA[33]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 137.345 76.575 137.545 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 137.345 76.575 137.545 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 137.345 76.575 137.545 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[33]

 PIN QA[34]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 140.795 76.575 140.995 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 140.795 76.575 140.995 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 140.795 76.575 140.995 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[34]

 PIN QA[35]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 141.885 76.575 142.085 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 141.885 76.575 142.085 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 141.885 76.575 142.085 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[35]

 PIN QA[36]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 145.335 76.575 145.535 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 145.335 76.575 145.535 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 145.335 76.575 145.535 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[36]

 PIN QA[37]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 146.425 76.575 146.625 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 146.425 76.575 146.625 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 146.425 76.575 146.625 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[37]

 PIN QA[38]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 149.875 76.575 150.075 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 149.875 76.575 150.075 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 149.875 76.575 150.075 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[38]

 PIN QA[39]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 150.965 76.575 151.165 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 150.965 76.575 151.165 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 150.965 76.575 151.165 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[39]

 PIN QA[40]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 154.415 76.575 154.615 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 154.415 76.575 154.615 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 154.415 76.575 154.615 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[40]

 PIN QA[41]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 155.505 76.575 155.705 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 155.505 76.575 155.705 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 155.505 76.575 155.705 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[41]

 PIN QA[42]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 158.955 76.575 159.155 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 158.955 76.575 159.155 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 158.955 76.575 159.155 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[42]

 PIN QA[43]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 160.045 76.575 160.245 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 160.045 76.575 160.245 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 160.045 76.575 160.245 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[43]

 PIN QA[44]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 163.495 76.575 163.695 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 163.495 76.575 163.695 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 163.495 76.575 163.695 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[44]

 PIN QA[45]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 164.585 76.575 164.785 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 164.585 76.575 164.785 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 164.585 76.575 164.785 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[45]

 PIN QA[46]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 168.035 76.575 168.235 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 168.035 76.575 168.235 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 168.035 76.575 168.235 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[46]

 PIN QA[47]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 169.125 76.575 169.325 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 169.125 76.575 169.325 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 169.125 76.575 169.325 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[47]

 PIN QA[48]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 172.575 76.575 172.775 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 172.575 76.575 172.775 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 172.575 76.575 172.775 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[48]

 PIN QA[49]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 173.665 76.575 173.865 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 173.665 76.575 173.865 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 173.665 76.575 173.865 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[49]

 PIN QA[50]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 177.115 76.575 177.315 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 177.115 76.575 177.315 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 177.115 76.575 177.315 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[50]

 PIN QA[51]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 178.205 76.575 178.405 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 178.205 76.575 178.405 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 178.205 76.575 178.405 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[51]

 PIN QA[52]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 181.655 76.575 181.855 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 181.655 76.575 181.855 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 181.655 76.575 181.855 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[52]

 PIN QA[53]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 182.745 76.575 182.945 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 182.745 76.575 182.945 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 182.745 76.575 182.945 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[53]

 PIN QA[54]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 186.195 76.575 186.395 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 186.195 76.575 186.395 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 186.195 76.575 186.395 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[54]

 PIN QA[55]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 187.285 76.575 187.485 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 187.285 76.575 187.485 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 187.285 76.575 187.485 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[55]

 PIN QA[56]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 190.735 76.575 190.935 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 190.735 76.575 190.935 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 190.735 76.575 190.935 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[56]

 PIN QA[57]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 191.825 76.575 192.025 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 191.825 76.575 192.025 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 191.825 76.575 192.025 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[57]

 PIN QA[58]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 195.275 76.575 195.475 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 195.275 76.575 195.475 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 195.275 76.575 195.475 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[58]

 PIN QA[59]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 196.365 76.575 196.565 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 196.365 76.575 196.565 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 196.365 76.575 196.565 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[59]

 PIN QA[60]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 199.815 76.575 200.015 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 199.815 76.575 200.015 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 199.815 76.575 200.015 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[60]

 PIN QA[61]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 200.905 76.575 201.105 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 200.905 76.575 201.105 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 200.905 76.575 201.105 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[61]

 PIN QA[62]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 204.355 76.575 204.555 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 204.355 76.575 204.555 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 204.355 76.575 204.555 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[62]

 PIN QA[63]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 205.445 76.575 205.645 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 205.445 76.575 205.645 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 205.445 76.575 205.645 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[63]

 PIN DB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[0]

 PIN DB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[1]

 PIN DB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[2]

 PIN DB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[3]

 PIN DB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[4]

 PIN DB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[5]

 PIN DB[6]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[6]

 PIN DB[7]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[7]

 PIN DB[8]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[8]

 PIN DB[9]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[9]

 PIN DB[10]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[10]

 PIN DB[11]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[11]

 PIN DB[12]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[12]

 PIN DB[13]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[13]

 PIN DB[14]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[14]

 PIN DB[15]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[15]

 PIN DB[16]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 40.13 0 40.33 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 40.13 0 40.33 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 40.13 0 40.33 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[16]

 PIN DB[17]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 41.71 0 41.91 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 41.71 0 41.91 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 41.71 0 41.91 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[17]

 PIN DB[18]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 44.67 0 44.87 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 44.67 0 44.87 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 44.67 0 44.87 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[18]

 PIN DB[19]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 46.25 0 46.45 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 46.25 0 46.45 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 46.25 0 46.45 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[19]

 PIN DB[20]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 49.21 0 49.41 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 49.21 0 49.41 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 49.21 0 49.41 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[20]

 PIN DB[21]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 50.79 0 50.99 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 50.79 0 50.99 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 50.79 0 50.99 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[21]

 PIN DB[22]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 53.75 0 53.95 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 53.75 0 53.95 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 53.75 0 53.95 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[22]

 PIN DB[23]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 55.33 0 55.53 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 55.33 0 55.53 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 55.33 0 55.53 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[23]

 PIN DB[24]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.29 0 58.49 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.29 0 58.49 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.29 0 58.49 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[24]

 PIN DB[25]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 59.87 0 60.07 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 59.87 0 60.07 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 59.87 0 60.07 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[25]

 PIN DB[26]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 62.83 0 63.03 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 62.83 0 63.03 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 62.83 0 63.03 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[26]

 PIN DB[27]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 64.41 0 64.61 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 64.41 0 64.61 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 64.41 0 64.61 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[27]

 PIN DB[28]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 67.37 0 67.57 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 67.37 0 67.57 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 67.37 0 67.57 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[28]

 PIN DB[29]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 68.95 0 69.15 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 68.95 0 69.15 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 68.95 0 69.15 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[29]

 PIN DB[30]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 71.91 0 72.11 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 71.91 0 72.11 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 71.91 0 72.11 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[30]

 PIN DB[31]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 73.49 0 73.69 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 73.49 0 73.69 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 73.49 0 73.69 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[31]

 PIN CLKB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 78.33 0 78.53 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 78.33 0 78.53 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 78.33 0 78.53 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKB

 PIN CENB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 78.82 0 79.02 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 78.82 0 79.02 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 78.82 0 79.02 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENB

 PIN AB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 100.43 0 100.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 100.43 0 100.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 100.43 0 100.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[5]

 PIN AB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 103.92 0 104.12 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 103.92 0 104.12 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 103.92 0 104.12 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[3]

 PIN AB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 105.355 0 105.555 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 105.355 0 105.555 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 105.355 0 105.555 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[4]

 PIN AB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 111.255 0 111.455 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 111.255 0 111.455 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 111.255 0 111.455 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[2]

 PIN AB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 111.905 0 112.105 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 111.905 0 112.105 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 111.905 0 112.105 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[0]

 PIN AB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 115.01 0 115.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 115.01 0 115.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 115.01 0 115.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[1]

 PIN DB[32]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 136.01 0 136.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 136.01 0 136.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 136.01 0 136.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[32]

 PIN DB[33]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 137.59 0 137.79 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 137.59 0 137.79 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 137.59 0 137.79 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[33]

 PIN DB[34]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 140.55 0 140.75 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 140.55 0 140.75 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 140.55 0 140.75 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[34]

 PIN DB[35]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 142.13 0 142.33 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 142.13 0 142.33 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 142.13 0 142.33 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[35]

 PIN DB[36]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 145.09 0 145.29 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 145.09 0 145.29 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 145.09 0 145.29 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[36]

 PIN DB[37]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 146.67 0 146.87 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 146.67 0 146.87 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 146.67 0 146.87 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[37]

 PIN DB[38]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 149.63 0 149.83 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 149.63 0 149.83 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 149.63 0 149.83 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[38]

 PIN DB[39]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 151.21 0 151.41 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 151.21 0 151.41 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 151.21 0 151.41 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[39]

 PIN DB[40]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 154.17 0 154.37 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 154.17 0 154.37 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 154.17 0 154.37 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[40]

 PIN DB[41]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 155.75 0 155.95 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 155.75 0 155.95 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 155.75 0 155.95 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[41]

 PIN DB[42]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 158.71 0 158.91 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 158.71 0 158.91 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 158.71 0 158.91 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[42]

 PIN DB[43]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 160.29 0 160.49 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 160.29 0 160.49 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 160.29 0 160.49 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[43]

 PIN DB[44]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 163.25 0 163.45 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 163.25 0 163.45 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 163.25 0 163.45 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[44]

 PIN DB[45]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 164.83 0 165.03 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 164.83 0 165.03 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 164.83 0 165.03 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[45]

 PIN DB[46]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 167.79 0 167.99 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 167.79 0 167.99 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 167.79 0 167.99 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[46]

 PIN DB[47]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 169.37 0 169.57 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 169.37 0 169.57 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 169.37 0 169.57 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[47]

 PIN DB[48]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 172.33 0 172.53 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 172.33 0 172.53 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 172.33 0 172.53 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[48]

 PIN DB[49]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 173.91 0 174.11 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 173.91 0 174.11 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 173.91 0 174.11 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[49]

 PIN DB[50]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 176.87 0 177.07 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 176.87 0 177.07 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 176.87 0 177.07 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[50]

 PIN DB[51]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 178.45 0 178.65 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 178.45 0 178.65 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 178.45 0 178.65 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[51]

 PIN DB[52]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 181.41 0 181.61 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 181.41 0 181.61 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 181.41 0 181.61 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[52]

 PIN DB[53]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 182.99 0 183.19 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 182.99 0 183.19 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 182.99 0 183.19 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[53]

 PIN DB[54]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 185.95 0 186.15 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 185.95 0 186.15 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 185.95 0 186.15 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[54]

 PIN DB[55]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 187.53 0 187.73 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 187.53 0 187.73 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 187.53 0 187.73 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[55]

 PIN DB[56]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 190.49 0 190.69 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 190.49 0 190.69 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 190.49 0 190.69 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[56]

 PIN DB[57]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 192.07 0 192.27 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 192.07 0 192.27 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 192.07 0 192.27 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[57]

 PIN DB[58]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 195.03 0 195.23 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 195.03 0 195.23 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 195.03 0 195.23 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[58]

 PIN DB[59]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 196.61 0 196.81 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 196.61 0 196.81 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 196.61 0 196.81 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[59]

 PIN DB[60]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 199.57 0 199.77 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 199.57 0 199.77 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 199.57 0 199.77 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[60]

 PIN DB[61]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 201.15 0 201.35 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 201.15 0 201.35 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 201.15 0 201.35 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[61]

 PIN DB[62]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 204.11 0 204.31 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 204.11 0 204.31 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 204.11 0 204.31 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[62]

 PIN DB[63]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 205.69 0 205.89 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 205.69 0 205.89 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 205.69 0 205.89 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[63]

 PIN VDD
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 2.43 0 3.93 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.01 0 11.51 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 11.51 0 13.01 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 19.09 0 20.59 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 20.59 0 22.09 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 28.17 0 29.67 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 29.67 0 31.17 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 37.25 0 38.75 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 38.75 0 40.25 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 46.33 0 47.83 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 47.83 0 49.33 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 55.41 0 56.91 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 56.91 0 58.41 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 64.49 0 65.99 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 65.99 0 67.49 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 73.57 0 75.07 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 78.29 0 83.29 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 88.74 0 92.24 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 96.44 0 100.44 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 109.26 0 113.26 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 117.46 0 120.96 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 126.41 0 131.41 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 134.63 0 136.13 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 142.21 0 143.71 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 143.71 0 145.21 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 151.29 0 152.79 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 152.79 0 154.29 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 160.37 0 161.87 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 161.87 0 163.37 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 169.45 0 170.95 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 170.95 0 172.45 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 178.53 0 180.03 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 180.03 0 181.53 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 187.61 0 189.11 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 189.11 0 190.61 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 196.69 0 198.19 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 198.19 0 199.69 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 205.77 0 207.27 76.575 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 5.47 0 6.97 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 6.97 0 8.47 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 14.55 0 16.05 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 16.05 0 17.55 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 23.63 0 25.13 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 25.13 0 26.63 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 32.71 0 34.21 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 34.21 0 35.71 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 41.79 0 43.29 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 43.29 0 44.79 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 50.87 0 52.37 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 52.37 0 53.87 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 59.95 0 61.45 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 61.45 0 62.95 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 69.03 0 70.53 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 70.53 0 72.03 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 84.14 0 88.14 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 92.84 0 95.84 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 101.845 0 107.845 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 113.86 0 116.86 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 121.56 0 125.56 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 137.67 0 139.17 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 139.17 0 140.67 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 146.75 0 148.25 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 148.25 0 149.75 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 155.83 0 157.33 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 157.33 0 158.83 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 164.91 0 166.41 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 166.41 0 167.91 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 173.99 0 175.49 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 175.49 0 176.99 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 183.07 0 184.57 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 184.57 0 186.07 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 192.15 0 193.65 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 193.65 0 195.15 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 201.23 0 202.73 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 202.73 0 204.23 76.575 ;      
 END
 END VSS

 OBS
 LAYER M1 ;
 RECT 0 0 3.72 0.585 ;
 RECT 4.1 0 5.3 0.585 ;
 RECT 5.68 0 8.26 0.585 ;
 RECT 8.64 0 9.84 0.585 ;
 RECT 10.22 0 12.8 0.585 ;
 RECT 13.18 0 14.38 0.585 ;
 RECT 14.76 0 17.34 0.585 ;
 RECT 17.72 0 18.92 0.585 ;
 RECT 19.3 0 21.88 0.585 ;
 RECT 22.26 0 23.46 0.585 ;
 RECT 23.84 0 26.42 0.585 ;
 RECT 26.8 0 28 0.585 ;
 RECT 28.38 0 30.96 0.585 ;
 RECT 31.34 0 32.54 0.585 ;
 RECT 32.92 0 35.5 0.585 ;
 RECT 35.88 0 37.08 0.585 ;
 RECT 37.46 0 40.04 0.585 ;
 RECT 40.42 0 41.62 0.585 ;
 RECT 42 0 44.58 0.585 ;
 RECT 44.96 0 46.16 0.585 ;
 RECT 46.54 0 49.12 0.585 ;
 RECT 49.5 0 50.7 0.585 ;
 RECT 51.08 0 53.66 0.585 ;
 RECT 54.04 0 55.24 0.585 ;
 RECT 55.62 0 58.2 0.585 ;
 RECT 58.58 0 59.78 0.585 ;
 RECT 60.16 0 62.74 0.585 ;
 RECT 63.12 0 64.32 0.585 ;
 RECT 64.7 0 67.28 0.585 ;
 RECT 67.66 0 68.86 0.585 ;
 RECT 69.24 0 71.82 0.585 ;
 RECT 72.2 0 73.4 0.585 ;
 RECT 73.78 0 78.24 0.585 ;
 RECT 78.62 0 78.73 0.585 ;
 RECT 79.11 0 100.34 0.585 ;
 RECT 100.72 0 103.83 0.585 ;
 RECT 104.21 0 105.265 0.585 ;
 RECT 105.645 0 111.165 0.585 ;
 RECT 111.545 0 111.815 0.585 ;
 RECT 112.195 0 114.92 0.585 ;
 RECT 115.3 0 135.92 0.585 ;
 RECT 136.3 0 137.5 0.585 ;
 RECT 137.88 0 140.46 0.585 ;
 RECT 140.84 0 142.04 0.585 ;
 RECT 142.42 0 145 0.585 ;
 RECT 145.38 0 146.58 0.585 ;
 RECT 146.96 0 149.54 0.585 ;
 RECT 149.92 0 151.12 0.585 ;
 RECT 151.5 0 154.08 0.585 ;
 RECT 154.46 0 155.66 0.585 ;
 RECT 156.04 0 158.62 0.585 ;
 RECT 159 0 160.2 0.585 ;
 RECT 160.58 0 163.16 0.585 ;
 RECT 163.54 0 164.74 0.585 ;
 RECT 165.12 0 167.7 0.585 ;
 RECT 168.08 0 169.28 0.585 ;
 RECT 169.66 0 172.24 0.585 ;
 RECT 172.62 0 173.82 0.585 ;
 RECT 174.2 0 176.78 0.585 ;
 RECT 177.16 0 178.36 0.585 ;
 RECT 178.74 0 181.32 0.585 ;
 RECT 181.7 0 182.9 0.585 ;
 RECT 183.28 0 185.86 0.585 ;
 RECT 186.24 0 187.44 0.585 ;
 RECT 187.82 0 190.4 0.585 ;
 RECT 190.78 0 191.98 0.585 ;
 RECT 192.36 0 194.94 0.585 ;
 RECT 195.32 0 196.52 0.585 ;
 RECT 196.9 0 199.48 0.585 ;
 RECT 199.86 0 201.06 0.585 ;
 RECT 201.44 0 204.02 0.585 ;
 RECT 204.4 0 205.6 0.585 ;
 RECT 205.98 0 209.7 0.585 ;
 RECT 0 76.575 3.965 75.99 ;
 RECT 4.345 76.575 5.055 75.99 ;
 RECT 5.435 76.575 8.505 75.99 ;
 RECT 8.885 76.575 9.595 75.99 ;
 RECT 9.975 76.575 13.045 75.99 ;
 RECT 13.425 76.575 14.135 75.99 ;
 RECT 14.515 76.575 17.585 75.99 ;
 RECT 17.965 76.575 18.675 75.99 ;
 RECT 19.055 76.575 22.125 75.99 ;
 RECT 22.505 76.575 23.215 75.99 ;
 RECT 23.595 76.575 26.665 75.99 ;
 RECT 27.045 76.575 27.755 75.99 ;
 RECT 28.135 76.575 31.205 75.99 ;
 RECT 31.585 76.575 32.295 75.99 ;
 RECT 32.675 76.575 35.745 75.99 ;
 RECT 36.125 76.575 36.835 75.99 ;
 RECT 37.215 76.575 40.285 75.99 ;
 RECT 40.665 76.575 41.375 75.99 ;
 RECT 41.755 76.575 44.825 75.99 ;
 RECT 45.205 76.575 45.915 75.99 ;
 RECT 46.295 76.575 49.365 75.99 ;
 RECT 49.745 76.575 50.455 75.99 ;
 RECT 50.835 76.575 53.905 75.99 ;
 RECT 54.285 76.575 54.995 75.99 ;
 RECT 55.375 76.575 58.445 75.99 ;
 RECT 58.825 76.575 59.535 75.99 ;
 RECT 59.915 76.575 62.985 75.99 ;
 RECT 63.365 76.575 64.075 75.99 ;
 RECT 64.455 76.575 67.525 75.99 ;
 RECT 67.905 76.575 68.615 75.99 ;
 RECT 68.995 76.575 72.065 75.99 ;
 RECT 72.445 76.575 73.155 75.99 ;
 RECT 73.535 76.575 91.445 75.99 ;
 RECT 91.825 76.575 94.55 75.99 ;
 RECT 94.93 76.575 95.2 75.99 ;
 RECT 95.58 76.575 101.1 75.99 ;
 RECT 101.48 76.575 102.535 75.99 ;
 RECT 102.915 76.575 106.025 75.99 ;
 RECT 106.405 76.575 127.86 75.99 ;
 RECT 128.24 76.575 128.35 75.99 ;
 RECT 128.73 76.575 136.165 75.99 ;
 RECT 136.545 76.575 137.255 75.99 ;
 RECT 137.635 76.575 140.705 75.99 ;
 RECT 141.085 76.575 141.795 75.99 ;
 RECT 142.175 76.575 145.245 75.99 ;
 RECT 145.625 76.575 146.335 75.99 ;
 RECT 146.715 76.575 149.785 75.99 ;
 RECT 150.165 76.575 150.875 75.99 ;
 RECT 151.255 76.575 154.325 75.99 ;
 RECT 154.705 76.575 155.415 75.99 ;
 RECT 155.795 76.575 158.865 75.99 ;
 RECT 159.245 76.575 159.955 75.99 ;
 RECT 160.335 76.575 163.405 75.99 ;
 RECT 163.785 76.575 164.495 75.99 ;
 RECT 164.875 76.575 167.945 75.99 ;
 RECT 168.325 76.575 169.035 75.99 ;
 RECT 169.415 76.575 172.485 75.99 ;
 RECT 172.865 76.575 173.575 75.99 ;
 RECT 173.955 76.575 177.025 75.99 ;
 RECT 177.405 76.575 178.115 75.99 ;
 RECT 178.495 76.575 181.565 75.99 ;
 RECT 181.945 76.575 182.655 75.99 ;
 RECT 183.035 76.575 186.105 75.99 ;
 RECT 186.485 76.575 187.195 75.99 ;
 RECT 187.575 76.575 190.645 75.99 ;
 RECT 191.025 76.575 191.735 75.99 ;
 RECT 192.115 76.575 195.185 75.99 ;
 RECT 195.565 76.575 196.275 75.99 ;
 RECT 196.655 76.575 199.725 75.99 ;
 RECT 200.105 76.575 200.815 75.99 ;
 RECT 201.195 76.575 204.265 75.99 ;
 RECT 204.645 76.575 205.355 75.99 ;
 RECT 205.735 76.575 209.7 75.99 ;
 RECT 0 0.585 209.7 75.99 ;
 LAYER M2 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 40.03 0.595 ;
 RECT 40.43 0 41.61 0.595 ;
 RECT 42.01 0 44.57 0.595 ;
 RECT 44.97 0 46.15 0.595 ;
 RECT 46.55 0 49.11 0.595 ;
 RECT 49.51 0 50.69 0.595 ;
 RECT 51.09 0 53.65 0.595 ;
 RECT 54.05 0 55.23 0.595 ;
 RECT 55.63 0 58.19 0.595 ;
 RECT 58.59 0 59.77 0.595 ;
 RECT 60.17 0 62.73 0.595 ;
 RECT 63.13 0 64.31 0.595 ;
 RECT 64.71 0 67.27 0.595 ;
 RECT 67.67 0 68.85 0.595 ;
 RECT 69.25 0 71.81 0.595 ;
 RECT 72.21 0 73.39 0.595 ;
 RECT 73.79 0 78.23 0.595 ;
 RECT 79.12 0 100.33 0.595 ;
 RECT 100.73 0 103.82 0.595 ;
 RECT 104.22 0 105.255 0.595 ;
 RECT 105.655 0 111.155 0.595 ;
 RECT 111.555 0 111.805 0.595 ;
 RECT 112.205 0 114.91 0.595 ;
 RECT 115.31 0 135.91 0.595 ;
 RECT 136.31 0 137.49 0.595 ;
 RECT 137.89 0 140.45 0.595 ;
 RECT 140.85 0 142.03 0.595 ;
 RECT 142.43 0 144.99 0.595 ;
 RECT 145.39 0 146.57 0.595 ;
 RECT 146.97 0 149.53 0.595 ;
 RECT 149.93 0 151.11 0.595 ;
 RECT 151.51 0 154.07 0.595 ;
 RECT 154.47 0 155.65 0.595 ;
 RECT 156.05 0 158.61 0.595 ;
 RECT 159.01 0 160.19 0.595 ;
 RECT 160.59 0 163.15 0.595 ;
 RECT 163.55 0 164.73 0.595 ;
 RECT 165.13 0 167.69 0.595 ;
 RECT 168.09 0 169.27 0.595 ;
 RECT 169.67 0 172.23 0.595 ;
 RECT 172.63 0 173.81 0.595 ;
 RECT 174.21 0 176.77 0.595 ;
 RECT 177.17 0 178.35 0.595 ;
 RECT 178.75 0 181.31 0.595 ;
 RECT 181.71 0 182.89 0.595 ;
 RECT 183.29 0 185.85 0.595 ;
 RECT 186.25 0 187.43 0.595 ;
 RECT 187.83 0 190.39 0.595 ;
 RECT 190.79 0 191.97 0.595 ;
 RECT 192.37 0 194.93 0.595 ;
 RECT 195.33 0 196.51 0.595 ;
 RECT 196.91 0 199.47 0.595 ;
 RECT 199.87 0 201.05 0.595 ;
 RECT 201.45 0 204.01 0.595 ;
 RECT 204.41 0 205.59 0.595 ;
 RECT 205.99 0 209.7 0.595 ;
 RECT 0 76.575 3.955 75.98 ;
 RECT 4.355 76.575 5.045 75.98 ;
 RECT 5.445 76.575 8.495 75.98 ;
 RECT 8.895 76.575 9.585 75.98 ;
 RECT 9.985 76.575 13.035 75.98 ;
 RECT 13.435 76.575 14.125 75.98 ;
 RECT 14.525 76.575 17.575 75.98 ;
 RECT 17.975 76.575 18.665 75.98 ;
 RECT 19.065 76.575 22.115 75.98 ;
 RECT 22.515 76.575 23.205 75.98 ;
 RECT 23.605 76.575 26.655 75.98 ;
 RECT 27.055 76.575 27.745 75.98 ;
 RECT 28.145 76.575 31.195 75.98 ;
 RECT 31.595 76.575 32.285 75.98 ;
 RECT 32.685 76.575 35.735 75.98 ;
 RECT 36.135 76.575 36.825 75.98 ;
 RECT 37.225 76.575 40.275 75.98 ;
 RECT 40.675 76.575 41.365 75.98 ;
 RECT 41.765 76.575 44.815 75.98 ;
 RECT 45.215 76.575 45.905 75.98 ;
 RECT 46.305 76.575 49.355 75.98 ;
 RECT 49.755 76.575 50.445 75.98 ;
 RECT 50.845 76.575 53.895 75.98 ;
 RECT 54.295 76.575 54.985 75.98 ;
 RECT 55.385 76.575 58.435 75.98 ;
 RECT 58.835 76.575 59.525 75.98 ;
 RECT 59.925 76.575 62.975 75.98 ;
 RECT 63.375 76.575 64.065 75.98 ;
 RECT 64.465 76.575 67.515 75.98 ;
 RECT 67.915 76.575 68.605 75.98 ;
 RECT 69.005 76.575 72.055 75.98 ;
 RECT 72.455 76.575 73.145 75.98 ;
 RECT 73.545 76.575 91.435 75.98 ;
 RECT 91.835 76.575 94.54 75.98 ;
 RECT 94.94 76.575 95.19 75.98 ;
 RECT 95.59 76.575 101.09 75.98 ;
 RECT 101.49 76.575 102.525 75.98 ;
 RECT 102.925 76.575 106.015 75.98 ;
 RECT 106.415 76.575 127.85 75.98 ;
 RECT 128.74 76.575 136.155 75.98 ;
 RECT 136.555 76.575 137.245 75.98 ;
 RECT 137.645 76.575 140.695 75.98 ;
 RECT 141.095 76.575 141.785 75.98 ;
 RECT 142.185 76.575 145.235 75.98 ;
 RECT 145.635 76.575 146.325 75.98 ;
 RECT 146.725 76.575 149.775 75.98 ;
 RECT 150.175 76.575 150.865 75.98 ;
 RECT 151.265 76.575 154.315 75.98 ;
 RECT 154.715 76.575 155.405 75.98 ;
 RECT 155.805 76.575 158.855 75.98 ;
 RECT 159.255 76.575 159.945 75.98 ;
 RECT 160.345 76.575 163.395 75.98 ;
 RECT 163.795 76.575 164.485 75.98 ;
 RECT 164.885 76.575 167.935 75.98 ;
 RECT 168.335 76.575 169.025 75.98 ;
 RECT 169.425 76.575 172.475 75.98 ;
 RECT 172.875 76.575 173.565 75.98 ;
 RECT 173.965 76.575 177.015 75.98 ;
 RECT 177.415 76.575 178.105 75.98 ;
 RECT 178.505 76.575 181.555 75.98 ;
 RECT 181.955 76.575 182.645 75.98 ;
 RECT 183.045 76.575 186.095 75.98 ;
 RECT 186.495 76.575 187.185 75.98 ;
 RECT 187.585 76.575 190.635 75.98 ;
 RECT 191.035 76.575 191.725 75.98 ;
 RECT 192.125 76.575 195.175 75.98 ;
 RECT 195.575 76.575 196.265 75.98 ;
 RECT 196.665 76.575 199.715 75.98 ;
 RECT 200.115 76.575 200.805 75.98 ;
 RECT 201.205 76.575 204.255 75.98 ;
 RECT 204.655 76.575 205.345 75.98 ;
 RECT 205.745 76.575 209.7 75.98 ;
 RECT 0 0.595 209.7 75.98 ;
 LAYER M3 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 40.03 0.595 ;
 RECT 40.43 0 41.61 0.595 ;
 RECT 42.01 0 44.57 0.595 ;
 RECT 44.97 0 46.15 0.595 ;
 RECT 46.55 0 49.11 0.595 ;
 RECT 49.51 0 50.69 0.595 ;
 RECT 51.09 0 53.65 0.595 ;
 RECT 54.05 0 55.23 0.595 ;
 RECT 55.63 0 58.19 0.595 ;
 RECT 58.59 0 59.77 0.595 ;
 RECT 60.17 0 62.73 0.595 ;
 RECT 63.13 0 64.31 0.595 ;
 RECT 64.71 0 67.27 0.595 ;
 RECT 67.67 0 68.85 0.595 ;
 RECT 69.25 0 71.81 0.595 ;
 RECT 72.21 0 73.39 0.595 ;
 RECT 73.79 0 78.23 0.595 ;
 RECT 79.12 0 100.33 0.595 ;
 RECT 100.73 0 103.82 0.595 ;
 RECT 104.22 0 105.255 0.595 ;
 RECT 105.655 0 111.155 0.595 ;
 RECT 111.555 0 111.805 0.595 ;
 RECT 112.205 0 114.91 0.595 ;
 RECT 115.31 0 135.91 0.595 ;
 RECT 136.31 0 137.49 0.595 ;
 RECT 137.89 0 140.45 0.595 ;
 RECT 140.85 0 142.03 0.595 ;
 RECT 142.43 0 144.99 0.595 ;
 RECT 145.39 0 146.57 0.595 ;
 RECT 146.97 0 149.53 0.595 ;
 RECT 149.93 0 151.11 0.595 ;
 RECT 151.51 0 154.07 0.595 ;
 RECT 154.47 0 155.65 0.595 ;
 RECT 156.05 0 158.61 0.595 ;
 RECT 159.01 0 160.19 0.595 ;
 RECT 160.59 0 163.15 0.595 ;
 RECT 163.55 0 164.73 0.595 ;
 RECT 165.13 0 167.69 0.595 ;
 RECT 168.09 0 169.27 0.595 ;
 RECT 169.67 0 172.23 0.595 ;
 RECT 172.63 0 173.81 0.595 ;
 RECT 174.21 0 176.77 0.595 ;
 RECT 177.17 0 178.35 0.595 ;
 RECT 178.75 0 181.31 0.595 ;
 RECT 181.71 0 182.89 0.595 ;
 RECT 183.29 0 185.85 0.595 ;
 RECT 186.25 0 187.43 0.595 ;
 RECT 187.83 0 190.39 0.595 ;
 RECT 190.79 0 191.97 0.595 ;
 RECT 192.37 0 194.93 0.595 ;
 RECT 195.33 0 196.51 0.595 ;
 RECT 196.91 0 199.47 0.595 ;
 RECT 199.87 0 201.05 0.595 ;
 RECT 201.45 0 204.01 0.595 ;
 RECT 204.41 0 205.59 0.595 ;
 RECT 205.99 0 209.7 0.595 ;
 RECT 0 76.575 3.955 75.98 ;
 RECT 4.355 76.575 5.045 75.98 ;
 RECT 5.445 76.575 8.495 75.98 ;
 RECT 8.895 76.575 9.585 75.98 ;
 RECT 9.985 76.575 13.035 75.98 ;
 RECT 13.435 76.575 14.125 75.98 ;
 RECT 14.525 76.575 17.575 75.98 ;
 RECT 17.975 76.575 18.665 75.98 ;
 RECT 19.065 76.575 22.115 75.98 ;
 RECT 22.515 76.575 23.205 75.98 ;
 RECT 23.605 76.575 26.655 75.98 ;
 RECT 27.055 76.575 27.745 75.98 ;
 RECT 28.145 76.575 31.195 75.98 ;
 RECT 31.595 76.575 32.285 75.98 ;
 RECT 32.685 76.575 35.735 75.98 ;
 RECT 36.135 76.575 36.825 75.98 ;
 RECT 37.225 76.575 40.275 75.98 ;
 RECT 40.675 76.575 41.365 75.98 ;
 RECT 41.765 76.575 44.815 75.98 ;
 RECT 45.215 76.575 45.905 75.98 ;
 RECT 46.305 76.575 49.355 75.98 ;
 RECT 49.755 76.575 50.445 75.98 ;
 RECT 50.845 76.575 53.895 75.98 ;
 RECT 54.295 76.575 54.985 75.98 ;
 RECT 55.385 76.575 58.435 75.98 ;
 RECT 58.835 76.575 59.525 75.98 ;
 RECT 59.925 76.575 62.975 75.98 ;
 RECT 63.375 76.575 64.065 75.98 ;
 RECT 64.465 76.575 67.515 75.98 ;
 RECT 67.915 76.575 68.605 75.98 ;
 RECT 69.005 76.575 72.055 75.98 ;
 RECT 72.455 76.575 73.145 75.98 ;
 RECT 73.545 76.575 91.435 75.98 ;
 RECT 91.835 76.575 94.54 75.98 ;
 RECT 94.94 76.575 95.19 75.98 ;
 RECT 95.59 76.575 101.09 75.98 ;
 RECT 101.49 76.575 102.525 75.98 ;
 RECT 102.925 76.575 106.015 75.98 ;
 RECT 106.415 76.575 127.85 75.98 ;
 RECT 128.74 76.575 136.155 75.98 ;
 RECT 136.555 76.575 137.245 75.98 ;
 RECT 137.645 76.575 140.695 75.98 ;
 RECT 141.095 76.575 141.785 75.98 ;
 RECT 142.185 76.575 145.235 75.98 ;
 RECT 145.635 76.575 146.325 75.98 ;
 RECT 146.725 76.575 149.775 75.98 ;
 RECT 150.175 76.575 150.865 75.98 ;
 RECT 151.265 76.575 154.315 75.98 ;
 RECT 154.715 76.575 155.405 75.98 ;
 RECT 155.805 76.575 158.855 75.98 ;
 RECT 159.255 76.575 159.945 75.98 ;
 RECT 160.345 76.575 163.395 75.98 ;
 RECT 163.795 76.575 164.485 75.98 ;
 RECT 164.885 76.575 167.935 75.98 ;
 RECT 168.335 76.575 169.025 75.98 ;
 RECT 169.425 76.575 172.475 75.98 ;
 RECT 172.875 76.575 173.565 75.98 ;
 RECT 173.965 76.575 177.015 75.98 ;
 RECT 177.415 76.575 178.105 75.98 ;
 RECT 178.505 76.575 181.555 75.98 ;
 RECT 181.955 76.575 182.645 75.98 ;
 RECT 183.045 76.575 186.095 75.98 ;
 RECT 186.495 76.575 187.185 75.98 ;
 RECT 187.585 76.575 190.635 75.98 ;
 RECT 191.035 76.575 191.725 75.98 ;
 RECT 192.125 76.575 195.175 75.98 ;
 RECT 195.575 76.575 196.265 75.98 ;
 RECT 196.665 76.575 199.715 75.98 ;
 RECT 200.115 76.575 200.805 75.98 ;
 RECT 201.205 76.575 204.255 75.98 ;
 RECT 204.655 76.575 205.345 75.98 ;
 RECT 205.745 76.575 209.7 75.98 ;
 RECT 0 0.595 209.7 75.98 ;

 LAYER V1 ;
 RECT 0 0 209.7 76.575 ;
 LAYER V2 ;
 RECT 0 0 209.7 76.575 ;
 LAYER V3 ;
 RECT 0 0 209.7 76.575 ;

 LAYER M4 ;
 RECT 75.17 0 78.19 0.595 ;
 RECT 75.17 0.595 78.19 76.575 ;
 RECT 83.39 0 84.04 0.595 ;
 RECT 83.39 0.595 84.04 76.575 ;
 RECT 88.24 0 88.64 0.595 ;
 RECT 88.24 0.595 88.64 76.575 ;
 RECT 92.34 0 92.74 0.595 ;
 RECT 92.34 0.595 92.74 76.575 ;
 RECT 95.94 0 96.34 0.595 ;
 RECT 95.94 0.595 96.34 76.575 ;
 RECT 100.54 0 101.745 0.595 ;
 RECT 100.54 0.595 101.745 76.575 ;
 RECT 107.945 0 109.16 0.595 ;
 RECT 107.945 0.595 109.16 76.575 ;
 RECT 113.36 0 113.76 0.595 ;
 RECT 113.36 0.595 113.76 76.575 ;
 RECT 116.96 0 117.36 0.595 ;
 RECT 116.96 0.595 117.36 76.575 ;
 RECT 121.06 0 121.46 0.595 ;
 RECT 121.06 0.595 121.46 76.575 ;
 RECT 125.66 0 126.31 0.595 ;
 RECT 125.66 0.595 126.31 76.575 ;
 RECT 131.51 0 134.53 0.595 ;
 RECT 131.51 0.595 134.53 76.575 ;
 LAYER V4 ;
 RECT 75.17 0 78.19 0.595 ;
 RECT 75.17 0.595 78.19 76.575 ;
 RECT 83.39 0 84.04 0.595 ;
 RECT 83.39 0.595 84.04 76.575 ;
 RECT 88.24 0 88.64 0.595 ;
 RECT 88.24 0.595 88.64 76.575 ;
 RECT 92.34 0 92.74 0.595 ;
 RECT 92.34 0.595 92.74 76.575 ;
 RECT 95.94 0 96.34 0.595 ;
 RECT 95.94 0.595 96.34 76.575 ;
 RECT 100.54 0 101.745 0.595 ;
 RECT 100.54 0.595 101.745 76.575 ;
 RECT 107.945 0 109.16 0.595 ;
 RECT 107.945 0.595 109.16 76.575 ;
 RECT 113.36 0 113.76 0.595 ;
 RECT 113.36 0.595 113.76 76.575 ;
 RECT 116.96 0 117.36 0.595 ;
 RECT 116.96 0.595 117.36 76.575 ;
 RECT 121.06 0 121.46 0.595 ;
 RECT 121.06 0.595 121.46 76.575 ;
 RECT 125.66 0 126.31 0.595 ;
 RECT 125.66 0.595 126.31 76.575 ;
 RECT 131.51 0 134.53 0.595 ;
 RECT 131.51 0.595 134.53 76.575 ;
 END

END qspi_data_info_64_mem
END LIBRARY