/*
     Copyright (c) 2018 SMIC             
     Filename:      qspi_data_info_32_mem.lef
     IP code:       S55NLLG2PH
     Version:       1.1.0
     CreateDate:    Oct 28, 2018        
                    
    LEF for General 2-PORT SRAM
    SMIC 55nm LL Logic Process

    Configuration: -instname qspi_data_info_32_mem -rows 64 -bits 32 -mux 1 
    Redundancy: Off
    Bit-Write: Off
*/

# DISCLAIMER                                                                      
#                                                                                   
#   SMIC hereby provides the quality information to you but makes no claims,      
# promises or guarantees about the accuracy, completeness, or adequacy of the     
# information herein. The information contained herein is provided on an "AS IS"  
# basis without any warranty, and SMIC assumes no obligation to provide support   
# of any kind or otherwise maintain the information.                                
#   SMIC disclaims any representation that the information does not infringe any  
# intellectual property rights or proprietary rights of any third parties. SMIC   
# makes no other warranty, whether express, implied or statutory as to any        
# matter whatsoever, including but not limited to the accuracy or sufficiency of  
# any information or the merchantability and fitness for a particular purpose.    
# Neither SMIC nor any of its representatives shall be liable for any cause of    
# action incurred to connect to this service.                                       
#                                                                                 
# STATEMENT OF USE AND CONFIDENTIALITY                                              
#                                                                                   
#   The following/attached material contains confidential and proprietary           
# information of SMIC. This material is based upon information which SMIC           
# considers reliable, but SMIC neither represents nor warrants that such          
# information is accurate or complete, and it must not be relied upon as such.    
# This information was prepared for informational purposes and is for the use     
# by SMIC's customer only. SMIC reserves the right to make changes in the           
# information at any time without notice.                                           
#   No part of this information may be reproduced, transmitted, transcribed,        
# stored in a retrieval system, or translated into any human or computer           
# language, in any form or by any means, electronic, mechanical, magnetic,          
# optical, chemical, manual, or otherwise, without the prior written consent of   
# SMIC. Any unauthorized use or disclosure of this material is strictly             
# prohibited and may be unlawful. By accepting this material, the receiving         
# party shall be deemed to have acknowledged, accepted, and agreed to be bound    
# by the foregoing limitations and restrictions. Thank you.                         
#                                                                                   

VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO qspi_data_info_32_mem
 CLASS BLOCK ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SIZE 137.06 BY 76.575 ;

 PIN QA[0]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 4.055 76.575 4.255 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[0]

 PIN QA[1]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.145 76.575 5.345 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[1]

 PIN QA[2]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.595 76.575 8.795 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[2]

 PIN QA[3]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.685 76.575 9.885 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[3]

 PIN QA[4]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 13.135 76.575 13.335 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[4]

 PIN QA[5]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.225 76.575 14.425 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[5]

 PIN QA[6]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.675 76.575 17.875 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[6]

 PIN QA[7]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 18.765 76.575 18.965 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[7]

 PIN QA[8]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 22.215 76.575 22.415 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[8]

 PIN QA[9]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.305 76.575 23.505 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[9]

 PIN QA[10]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.755 76.575 26.955 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[10]

 PIN QA[11]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 27.845 76.575 28.045 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[11]

 PIN QA[12]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.295 76.575 31.495 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[12]

 PIN QA[13]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.385 76.575 32.585 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[13]

 PIN QA[14]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.835 76.575 36.035 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[14]

 PIN QA[15]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 36.925 76.575 37.125 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[15]

 PIN AA[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 55.215 76.575 55.415 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 55.215 76.575 55.415 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 55.215 76.575 55.415 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[1]

 PIN AA[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.32 76.575 58.52 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.32 76.575 58.52 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.32 76.575 58.52 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[0]

 PIN AA[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 58.97 76.575 59.17 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 58.97 76.575 59.17 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 58.97 76.575 59.17 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[2]

 PIN AA[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 64.87 76.575 65.07 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 64.87 76.575 65.07 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 64.87 76.575 65.07 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[4]

 PIN AA[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 66.305 76.575 66.505 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 66.305 76.575 66.505 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 66.305 76.575 66.505 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[3]

 PIN AA[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 69.795 76.575 69.995 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 69.795 76.575 69.995 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 69.795 76.575 69.995 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AA[5]

 PIN CENA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 91.63 76.575 91.83 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 91.63 76.575 91.83 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 91.63 76.575 91.83 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENA

 PIN CLKA
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 92.12 76.575 92.32 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 92.12 76.575 92.32 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 92.12 76.575 92.32 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKA

 PIN QA[16]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 99.935 76.575 100.135 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 99.935 76.575 100.135 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 99.935 76.575 100.135 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[16]

 PIN QA[17]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 101.025 76.575 101.225 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 101.025 76.575 101.225 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 101.025 76.575 101.225 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[17]

 PIN QA[18]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 104.475 76.575 104.675 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 104.475 76.575 104.675 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 104.475 76.575 104.675 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[18]

 PIN QA[19]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 105.565 76.575 105.765 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 105.565 76.575 105.765 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 105.565 76.575 105.765 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[19]

 PIN QA[20]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 109.015 76.575 109.215 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 109.015 76.575 109.215 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 109.015 76.575 109.215 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[20]

 PIN QA[21]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 110.105 76.575 110.305 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 110.105 76.575 110.305 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 110.105 76.575 110.305 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[21]

 PIN QA[22]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 113.555 76.575 113.755 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 113.555 76.575 113.755 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 113.555 76.575 113.755 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[22]

 PIN QA[23]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 114.645 76.575 114.845 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 114.645 76.575 114.845 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 114.645 76.575 114.845 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[23]

 PIN QA[24]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 118.095 76.575 118.295 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 118.095 76.575 118.295 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 118.095 76.575 118.295 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[24]

 PIN QA[25]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 119.185 76.575 119.385 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 119.185 76.575 119.385 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 119.185 76.575 119.385 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[25]

 PIN QA[26]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 122.635 76.575 122.835 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 122.635 76.575 122.835 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 122.635 76.575 122.835 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[26]

 PIN QA[27]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 123.725 76.575 123.925 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 123.725 76.575 123.925 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 123.725 76.575 123.925 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[27]

 PIN QA[28]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 127.175 76.575 127.375 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 127.175 76.575 127.375 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 127.175 76.575 127.375 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[28]

 PIN QA[29]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 128.265 76.575 128.465 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 128.265 76.575 128.465 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 128.265 76.575 128.465 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[29]

 PIN QA[30]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 131.715 76.575 131.915 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 131.715 76.575 131.915 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 131.715 76.575 131.915 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[30]

 PIN QA[31]
 DIRECTION OUTPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 132.805 76.575 133.005 76.08 ;
 END
 PORT
 LAYER M2 ;
 RECT 132.805 76.575 133.005 76.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 132.805 76.575 133.005 76.08 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END QA[31]

 PIN DB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 3.81 0 4.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[0]

 PIN DB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 5.39 0 5.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[1]

 PIN DB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 8.35 0 8.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[2]

 PIN DB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 9.93 0 10.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[3]

 PIN DB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 12.89 0 13.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[4]

 PIN DB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 14.47 0 14.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[5]

 PIN DB[6]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 17.43 0 17.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[6]

 PIN DB[7]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 19.01 0 19.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[7]

 PIN DB[8]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 21.97 0 22.17 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[8]

 PIN DB[9]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 23.55 0 23.75 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[9]

 PIN DB[10]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 26.51 0 26.71 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[10]

 PIN DB[11]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 28.09 0 28.29 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[11]

 PIN DB[12]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 31.05 0 31.25 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[12]

 PIN DB[13]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 32.63 0 32.83 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[13]

 PIN DB[14]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 35.59 0 35.79 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[14]

 PIN DB[15]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 37.17 0 37.37 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[15]

 PIN CLKB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.01 0 42.21 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CLKB

 PIN CENB
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 42.5 0 42.7 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END CENB

 PIN AB[5]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 64.11 0 64.31 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 64.11 0 64.31 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 64.11 0 64.31 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[5]

 PIN AB[3]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 67.6 0 67.8 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[3]

 PIN AB[4]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 69.035 0 69.235 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[4]

 PIN AB[2]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 74.935 0 75.135 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[2]

 PIN AB[0]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 75.585 0 75.785 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[0]

 PIN AB[1]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 78.69 0 78.89 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END AB[1]

 PIN DB[16]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 99.69 0 99.89 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[16]

 PIN DB[17]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 101.27 0 101.47 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[17]

 PIN DB[18]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 104.23 0 104.43 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[18]

 PIN DB[19]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 105.81 0 106.01 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[19]

 PIN DB[20]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 108.77 0 108.97 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[20]

 PIN DB[21]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 110.35 0 110.55 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[21]

 PIN DB[22]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 113.31 0 113.51 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[22]

 PIN DB[23]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 114.89 0 115.09 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[23]

 PIN DB[24]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 117.85 0 118.05 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[24]

 PIN DB[25]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 119.43 0 119.63 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[25]

 PIN DB[26]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 122.39 0 122.59 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[26]

 PIN DB[27]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 123.97 0 124.17 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[27]

 PIN DB[28]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 126.93 0 127.13 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[28]

 PIN DB[29]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 128.51 0 128.71 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[29]

 PIN DB[30]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 131.47 0 131.67 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[30]

 PIN DB[31]
 DIRECTION INPUT ;
 USE SIGNAL ; 
 PORT
 LAYER M3 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 PORT
 LAYER M2 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 PORT
 LAYER M1 ;
 RECT 133.05 0 133.25 0.495 ;
 END
 ANTENNAGATEAREA 0.025 ;
 ANTENNADIFFAREA 0.060 ; 
 END DB[31]

 PIN VDD
 USE POWER ;
 PORT
 LAYER M4 ;
 RECT 2.43 0 3.93 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 10.01 0 11.51 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 11.51 0 13.01 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 19.09 0 20.59 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 20.59 0 22.09 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 28.17 0 29.67 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 29.67 0 31.17 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 37.25 0 38.75 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 41.97 0 46.97 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 52.42 0 55.92 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 60.12 0 64.12 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 72.94 0 76.94 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 81.14 0 84.64 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 90.09 0 95.09 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 98.31 0 99.81 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 105.89 0 107.39 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 107.39 0 108.89 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 114.97 0 116.47 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 116.47 0 117.97 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 124.05 0 125.55 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 125.55 0 127.05 76.575 ;    
 END 
 PORT
 LAYER M4 ;
 RECT 133.13 0 134.63 76.575 ;    
 END 
 END VDD

 PIN VSS
 USE GROUND ;
 PORT
 LAYER M4 ;
 RECT 5.47 0 6.97 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 6.97 0 8.47 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 14.55 0 16.05 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 16.05 0 17.55 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 23.63 0 25.13 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 25.13 0 26.63 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 32.71 0 34.21 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 34.21 0 35.71 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 47.82 0 51.82 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 56.52 0 59.52 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 65.525 0 71.525 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 77.54 0 80.54 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 85.24 0 89.24 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 101.35 0 102.85 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 102.85 0 104.35 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 110.43 0 111.93 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 111.93 0 113.43 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 119.51 0 121.01 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 121.01 0 122.51 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 128.59 0 130.09 76.575 ;      
 END
 PORT
 LAYER M4 ;
 RECT 130.09 0 131.59 76.575 ;      
 END
 END VSS

 OBS
 LAYER M1 ;
 RECT 0 0 3.72 0.585 ;
 RECT 4.1 0 5.3 0.585 ;
 RECT 5.68 0 8.26 0.585 ;
 RECT 8.64 0 9.84 0.585 ;
 RECT 10.22 0 12.8 0.585 ;
 RECT 13.18 0 14.38 0.585 ;
 RECT 14.76 0 17.34 0.585 ;
 RECT 17.72 0 18.92 0.585 ;
 RECT 19.3 0 21.88 0.585 ;
 RECT 22.26 0 23.46 0.585 ;
 RECT 23.84 0 26.42 0.585 ;
 RECT 26.8 0 28 0.585 ;
 RECT 28.38 0 30.96 0.585 ;
 RECT 31.34 0 32.54 0.585 ;
 RECT 32.92 0 35.5 0.585 ;
 RECT 35.88 0 37.08 0.585 ;
 RECT 37.46 0 41.92 0.585 ;
 RECT 42.3 0 42.41 0.585 ;
 RECT 42.79 0 64.02 0.585 ;
 RECT 64.4 0 67.51 0.585 ;
 RECT 67.89 0 68.945 0.585 ;
 RECT 69.325 0 74.845 0.585 ;
 RECT 75.225 0 75.495 0.585 ;
 RECT 75.875 0 78.6 0.585 ;
 RECT 78.98 0 99.6 0.585 ;
 RECT 99.98 0 101.18 0.585 ;
 RECT 101.56 0 104.14 0.585 ;
 RECT 104.52 0 105.72 0.585 ;
 RECT 106.1 0 108.68 0.585 ;
 RECT 109.06 0 110.26 0.585 ;
 RECT 110.64 0 113.22 0.585 ;
 RECT 113.6 0 114.8 0.585 ;
 RECT 115.18 0 117.76 0.585 ;
 RECT 118.14 0 119.34 0.585 ;
 RECT 119.72 0 122.3 0.585 ;
 RECT 122.68 0 123.88 0.585 ;
 RECT 124.26 0 126.84 0.585 ;
 RECT 127.22 0 128.42 0.585 ;
 RECT 128.8 0 131.38 0.585 ;
 RECT 131.76 0 132.96 0.585 ;
 RECT 133.34 0 137.06 0.585 ;
 RECT 0 76.575 3.965 75.99 ;
 RECT 4.345 76.575 5.055 75.99 ;
 RECT 5.435 76.575 8.505 75.99 ;
 RECT 8.885 76.575 9.595 75.99 ;
 RECT 9.975 76.575 13.045 75.99 ;
 RECT 13.425 76.575 14.135 75.99 ;
 RECT 14.515 76.575 17.585 75.99 ;
 RECT 17.965 76.575 18.675 75.99 ;
 RECT 19.055 76.575 22.125 75.99 ;
 RECT 22.505 76.575 23.215 75.99 ;
 RECT 23.595 76.575 26.665 75.99 ;
 RECT 27.045 76.575 27.755 75.99 ;
 RECT 28.135 76.575 31.205 75.99 ;
 RECT 31.585 76.575 32.295 75.99 ;
 RECT 32.675 76.575 35.745 75.99 ;
 RECT 36.125 76.575 36.835 75.99 ;
 RECT 37.215 76.575 55.125 75.99 ;
 RECT 55.505 76.575 58.23 75.99 ;
 RECT 58.61 76.575 58.88 75.99 ;
 RECT 59.26 76.575 64.78 75.99 ;
 RECT 65.16 76.575 66.215 75.99 ;
 RECT 66.595 76.575 69.705 75.99 ;
 RECT 70.085 76.575 91.54 75.99 ;
 RECT 91.92 76.575 92.03 75.99 ;
 RECT 92.41 76.575 99.845 75.99 ;
 RECT 100.225 76.575 100.935 75.99 ;
 RECT 101.315 76.575 104.385 75.99 ;
 RECT 104.765 76.575 105.475 75.99 ;
 RECT 105.855 76.575 108.925 75.99 ;
 RECT 109.305 76.575 110.015 75.99 ;
 RECT 110.395 76.575 113.465 75.99 ;
 RECT 113.845 76.575 114.555 75.99 ;
 RECT 114.935 76.575 118.005 75.99 ;
 RECT 118.385 76.575 119.095 75.99 ;
 RECT 119.475 76.575 122.545 75.99 ;
 RECT 122.925 76.575 123.635 75.99 ;
 RECT 124.015 76.575 127.085 75.99 ;
 RECT 127.465 76.575 128.175 75.99 ;
 RECT 128.555 76.575 131.625 75.99 ;
 RECT 132.005 76.575 132.715 75.99 ;
 RECT 133.095 76.575 137.06 75.99 ;
 RECT 0 0.585 137.06 75.99 ;
 LAYER M2 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 41.91 0.595 ;
 RECT 42.8 0 64.01 0.595 ;
 RECT 64.41 0 67.5 0.595 ;
 RECT 67.9 0 68.935 0.595 ;
 RECT 69.335 0 74.835 0.595 ;
 RECT 75.235 0 75.485 0.595 ;
 RECT 75.885 0 78.59 0.595 ;
 RECT 78.99 0 99.59 0.595 ;
 RECT 99.99 0 101.17 0.595 ;
 RECT 101.57 0 104.13 0.595 ;
 RECT 104.53 0 105.71 0.595 ;
 RECT 106.11 0 108.67 0.595 ;
 RECT 109.07 0 110.25 0.595 ;
 RECT 110.65 0 113.21 0.595 ;
 RECT 113.61 0 114.79 0.595 ;
 RECT 115.19 0 117.75 0.595 ;
 RECT 118.15 0 119.33 0.595 ;
 RECT 119.73 0 122.29 0.595 ;
 RECT 122.69 0 123.87 0.595 ;
 RECT 124.27 0 126.83 0.595 ;
 RECT 127.23 0 128.41 0.595 ;
 RECT 128.81 0 131.37 0.595 ;
 RECT 131.77 0 132.95 0.595 ;
 RECT 133.35 0 137.06 0.595 ;
 RECT 0 76.575 3.955 75.98 ;
 RECT 4.355 76.575 5.045 75.98 ;
 RECT 5.445 76.575 8.495 75.98 ;
 RECT 8.895 76.575 9.585 75.98 ;
 RECT 9.985 76.575 13.035 75.98 ;
 RECT 13.435 76.575 14.125 75.98 ;
 RECT 14.525 76.575 17.575 75.98 ;
 RECT 17.975 76.575 18.665 75.98 ;
 RECT 19.065 76.575 22.115 75.98 ;
 RECT 22.515 76.575 23.205 75.98 ;
 RECT 23.605 76.575 26.655 75.98 ;
 RECT 27.055 76.575 27.745 75.98 ;
 RECT 28.145 76.575 31.195 75.98 ;
 RECT 31.595 76.575 32.285 75.98 ;
 RECT 32.685 76.575 35.735 75.98 ;
 RECT 36.135 76.575 36.825 75.98 ;
 RECT 37.225 76.575 55.115 75.98 ;
 RECT 55.515 76.575 58.22 75.98 ;
 RECT 58.62 76.575 58.87 75.98 ;
 RECT 59.27 76.575 64.77 75.98 ;
 RECT 65.17 76.575 66.205 75.98 ;
 RECT 66.605 76.575 69.695 75.98 ;
 RECT 70.095 76.575 91.53 75.98 ;
 RECT 92.42 76.575 99.835 75.98 ;
 RECT 100.235 76.575 100.925 75.98 ;
 RECT 101.325 76.575 104.375 75.98 ;
 RECT 104.775 76.575 105.465 75.98 ;
 RECT 105.865 76.575 108.915 75.98 ;
 RECT 109.315 76.575 110.005 75.98 ;
 RECT 110.405 76.575 113.455 75.98 ;
 RECT 113.855 76.575 114.545 75.98 ;
 RECT 114.945 76.575 117.995 75.98 ;
 RECT 118.395 76.575 119.085 75.98 ;
 RECT 119.485 76.575 122.535 75.98 ;
 RECT 122.935 76.575 123.625 75.98 ;
 RECT 124.025 76.575 127.075 75.98 ;
 RECT 127.475 76.575 128.165 75.98 ;
 RECT 128.565 76.575 131.615 75.98 ;
 RECT 132.015 76.575 132.705 75.98 ;
 RECT 133.105 76.575 137.06 75.98 ;
 RECT 0 0.595 137.06 75.98 ;
 LAYER M3 ;
 RECT 0 0 3.71 0.595 ;
 RECT 4.11 0 5.29 0.595 ;
 RECT 5.69 0 8.25 0.595 ;
 RECT 8.65 0 9.83 0.595 ;
 RECT 10.23 0 12.79 0.595 ;
 RECT 13.19 0 14.37 0.595 ;
 RECT 14.77 0 17.33 0.595 ;
 RECT 17.73 0 18.91 0.595 ;
 RECT 19.31 0 21.87 0.595 ;
 RECT 22.27 0 23.45 0.595 ;
 RECT 23.85 0 26.41 0.595 ;
 RECT 26.81 0 27.99 0.595 ;
 RECT 28.39 0 30.95 0.595 ;
 RECT 31.35 0 32.53 0.595 ;
 RECT 32.93 0 35.49 0.595 ;
 RECT 35.89 0 37.07 0.595 ;
 RECT 37.47 0 41.91 0.595 ;
 RECT 42.8 0 64.01 0.595 ;
 RECT 64.41 0 67.5 0.595 ;
 RECT 67.9 0 68.935 0.595 ;
 RECT 69.335 0 74.835 0.595 ;
 RECT 75.235 0 75.485 0.595 ;
 RECT 75.885 0 78.59 0.595 ;
 RECT 78.99 0 99.59 0.595 ;
 RECT 99.99 0 101.17 0.595 ;
 RECT 101.57 0 104.13 0.595 ;
 RECT 104.53 0 105.71 0.595 ;
 RECT 106.11 0 108.67 0.595 ;
 RECT 109.07 0 110.25 0.595 ;
 RECT 110.65 0 113.21 0.595 ;
 RECT 113.61 0 114.79 0.595 ;
 RECT 115.19 0 117.75 0.595 ;
 RECT 118.15 0 119.33 0.595 ;
 RECT 119.73 0 122.29 0.595 ;
 RECT 122.69 0 123.87 0.595 ;
 RECT 124.27 0 126.83 0.595 ;
 RECT 127.23 0 128.41 0.595 ;
 RECT 128.81 0 131.37 0.595 ;
 RECT 131.77 0 132.95 0.595 ;
 RECT 133.35 0 137.06 0.595 ;
 RECT 0 76.575 3.955 75.98 ;
 RECT 4.355 76.575 5.045 75.98 ;
 RECT 5.445 76.575 8.495 75.98 ;
 RECT 8.895 76.575 9.585 75.98 ;
 RECT 9.985 76.575 13.035 75.98 ;
 RECT 13.435 76.575 14.125 75.98 ;
 RECT 14.525 76.575 17.575 75.98 ;
 RECT 17.975 76.575 18.665 75.98 ;
 RECT 19.065 76.575 22.115 75.98 ;
 RECT 22.515 76.575 23.205 75.98 ;
 RECT 23.605 76.575 26.655 75.98 ;
 RECT 27.055 76.575 27.745 75.98 ;
 RECT 28.145 76.575 31.195 75.98 ;
 RECT 31.595 76.575 32.285 75.98 ;
 RECT 32.685 76.575 35.735 75.98 ;
 RECT 36.135 76.575 36.825 75.98 ;
 RECT 37.225 76.575 55.115 75.98 ;
 RECT 55.515 76.575 58.22 75.98 ;
 RECT 58.62 76.575 58.87 75.98 ;
 RECT 59.27 76.575 64.77 75.98 ;
 RECT 65.17 76.575 66.205 75.98 ;
 RECT 66.605 76.575 69.695 75.98 ;
 RECT 70.095 76.575 91.53 75.98 ;
 RECT 92.42 76.575 99.835 75.98 ;
 RECT 100.235 76.575 100.925 75.98 ;
 RECT 101.325 76.575 104.375 75.98 ;
 RECT 104.775 76.575 105.465 75.98 ;
 RECT 105.865 76.575 108.915 75.98 ;
 RECT 109.315 76.575 110.005 75.98 ;
 RECT 110.405 76.575 113.455 75.98 ;
 RECT 113.855 76.575 114.545 75.98 ;
 RECT 114.945 76.575 117.995 75.98 ;
 RECT 118.395 76.575 119.085 75.98 ;
 RECT 119.485 76.575 122.535 75.98 ;
 RECT 122.935 76.575 123.625 75.98 ;
 RECT 124.025 76.575 127.075 75.98 ;
 RECT 127.475 76.575 128.165 75.98 ;
 RECT 128.565 76.575 131.615 75.98 ;
 RECT 132.015 76.575 132.705 75.98 ;
 RECT 133.105 76.575 137.06 75.98 ;
 RECT 0 0.595 137.06 75.98 ;

 LAYER V1 ;
 RECT 0 0 137.06 76.575 ;
 LAYER V2 ;
 RECT 0 0 137.06 76.575 ;
 LAYER V3 ;
 RECT 0 0 137.06 76.575 ;

 LAYER M4 ;
 RECT 38.85 0 41.87 0.595 ;
 RECT 38.85 0.595 41.87 76.575 ;
 RECT 47.07 0 47.72 0.595 ;
 RECT 47.07 0.595 47.72 76.575 ;
 RECT 51.92 0 52.32 0.595 ;
 RECT 51.92 0.595 52.32 76.575 ;
 RECT 56.02 0 56.42 0.595 ;
 RECT 56.02 0.595 56.42 76.575 ;
 RECT 59.62 0 60.02 0.595 ;
 RECT 59.62 0.595 60.02 76.575 ;
 RECT 64.22 0 65.425 0.595 ;
 RECT 64.22 0.595 65.425 76.575 ;
 RECT 71.625 0 72.84 0.595 ;
 RECT 71.625 0.595 72.84 76.575 ;
 RECT 77.04 0 77.44 0.595 ;
 RECT 77.04 0.595 77.44 76.575 ;
 RECT 80.64 0 81.04 0.595 ;
 RECT 80.64 0.595 81.04 76.575 ;
 RECT 84.74 0 85.14 0.595 ;
 RECT 84.74 0.595 85.14 76.575 ;
 RECT 89.34 0 89.99 0.595 ;
 RECT 89.34 0.595 89.99 76.575 ;
 RECT 95.19 0 98.21 0.595 ;
 RECT 95.19 0.595 98.21 76.575 ;
 LAYER V4 ;
 RECT 38.85 0 41.87 0.595 ;
 RECT 38.85 0.595 41.87 76.575 ;
 RECT 47.07 0 47.72 0.595 ;
 RECT 47.07 0.595 47.72 76.575 ;
 RECT 51.92 0 52.32 0.595 ;
 RECT 51.92 0.595 52.32 76.575 ;
 RECT 56.02 0 56.42 0.595 ;
 RECT 56.02 0.595 56.42 76.575 ;
 RECT 59.62 0 60.02 0.595 ;
 RECT 59.62 0.595 60.02 76.575 ;
 RECT 64.22 0 65.425 0.595 ;
 RECT 64.22 0.595 65.425 76.575 ;
 RECT 71.625 0 72.84 0.595 ;
 RECT 71.625 0.595 72.84 76.575 ;
 RECT 77.04 0 77.44 0.595 ;
 RECT 77.04 0.595 77.44 76.575 ;
 RECT 80.64 0 81.04 0.595 ;
 RECT 80.64 0.595 81.04 76.575 ;
 RECT 84.74 0 85.14 0.595 ;
 RECT 84.74 0.595 85.14 76.575 ;
 RECT 89.34 0 89.99 0.595 ;
 RECT 89.34 0.595 89.99 76.575 ;
 RECT 95.19 0 98.21 0.595 ;
 RECT 95.19 0.595 98.21 76.575 ;
 END

END qspi_data_info_32_mem
END LIBRARY