*****************************************************************************
* CDL NETLIST:
* CELL NAME: qspi_data_info_32_mem
* IP code : S55NLLG2PH
*****************************************************************************


*****************************************************************************
* GLOBAL NET DECLARATIONS
*****************************************************************************


*****************************************************************************
* PIN CONTROL STATEMENT
*****************************************************************************


*****************************************************************************
* BIPOLAR DECLARATIONS
*****************************************************************************


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* Block: qspi_data_info_32_mem_TIE_LOW_X1                                          *
*******************************************************************************
.SUBCKT qspi_data_info_32_mem_TIE_LOW_X1 PULL0 VSS VDD
MP18 VDD NET2 NET2 VDD P12LL W=1.0U L=0.06U M=1
MN18 PULL0 NET2 VSS VSS N12LL W=1.5U L=0.06U M=1
.ENDS qspi_data_info_32_mem_TIE_LOW_X1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* Block: qspi_data_info_32_mem_TIE_HIGH_X1                                        *
*******************************************************************************
.SUBCKT qspi_data_info_32_mem_TIE_HIGH_X1 PULL1 VSS VDD
MP18 VDD NET2 PULL1 VDD P12LL W=2.0U L=0.06U M=1
MN18 NET2 NET2 VSS VSS N12LL W=1.0U L=0.06U M=1
.ENDS qspi_data_info_32_mem_TIE_HIGH_X1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* Block: qspi_data_info_32_mem_TIE_LOW_X2                                          *
*******************************************************************************
.SUBCKT qspi_data_info_32_mem_TIE_LOW_X2 PULL0 VSS VDD
MP18 VDD NET2 NET2 VDD P12LL W=0.4U L=0.06U M=1
MN18 PULL0 NET2 VSS VSS N12LL W=1U L=0.06U M=1
.ENDS qspi_data_info_32_mem_TIE_LOW_X2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_DISCHARGECELLS                                                    *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_DISCHARGECELLS VDD VSS DUM_BL EMCLK S[5] S[4] S[3] S[2] S[1] S[0]

M0 3 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=575 $Y=-500 $D=24
M1 3 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=575 $Y=1010 $D=24
M2 DUM_BL EMCLK 3 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=1795 $Y=-500 $D=24
M3 DUM_BL EMCLK 3 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=1795 $Y=1010 $D=24
M4 5 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=3345 $Y=-500 $D=24
M5 5 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=3345 $Y=1010 $D=24
M6 DUM_BL EMCLK 5 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=4565 $Y=-500 $D=24
M7 DUM_BL EMCLK 5 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=4565 $Y=1010 $D=24
M8 7 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=5855 $Y=-500 $D=24
M9 7 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=5855 $Y=1010 $D=24
M10 DUM_BL EMCLK 7 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=7075 $Y=-500 $D=24
M11 DUM_BL EMCLK 7 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=7075 $Y=1010 $D=24
M12 9 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=8625 $Y=-500 $D=24
M13 9 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=8625 $Y=1010 $D=24
M14 DUM_BL EMCLK 9 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=9845 $Y=-500 $D=24
M15 DUM_BL EMCLK 9 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=9845 $Y=1010 $D=24
M16 9 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=11150 $Y=-500 $D=24
M17 9 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=11150 $Y=1010 $D=24
M18 DUM_BL EMCLK 9 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=12370 $Y=-500 $D=24
M19 DUM_BL EMCLK 9 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=12370 $Y=1010 $D=24
M20 11 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=13920 $Y=-500 $D=24
M21 11 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=13920 $Y=1010 $D=24
M22 DUM_BL EMCLK 11 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=15140 $Y=-500 $D=24
M23 DUM_BL EMCLK 11 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=15140 $Y=1010 $D=24
M24 11 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=16430 $Y=-500 $D=24
M25 11 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=16430 $Y=1010 $D=24
M26 DUM_BL EMCLK 11 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=17650 $Y=-500 $D=24
M27 DUM_BL EMCLK 11 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=17650 $Y=1010 $D=24
M28 13 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=19200 $Y=-500 $D=24
M29 13 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=19200 $Y=1010 $D=24
M30 DUM_BL EMCLK 13 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=20420 $Y=-500 $D=24
M31 DUM_BL EMCLK 13 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=20420 $Y=1010 $D=24
M32 13 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=21795 $Y=-500 $D=24
M33 13 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=21795 $Y=1010 $D=24
M34 DUM_BL EMCLK 13 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=23015 $Y=-500 $D=24
M35 DUM_BL EMCLK 13 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=23015 $Y=1010 $D=24
M36 16 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=24565 $Y=-500 $D=24
M37 16 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=24565 $Y=1010 $D=24
M38 DUM_BL EMCLK 16 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=25785 $Y=-500 $D=24
M39 DUM_BL EMCLK 16 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=25785 $Y=1010 $D=24
M40 16 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=27075 $Y=-500 $D=24
M41 16 EMCLK DUM_BL VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=27075 $Y=1010 $D=24
M42 DUM_BL EMCLK 16 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=28295 $Y=-500 $D=24
M43 DUM_BL EMCLK 16 VSS RFNPGBHVT L=9E-08 W=1.2E-07 $X=28295 $Y=1010 $D=24
M44 VSS VDD 3 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=980 $Y=-840 $D=26
M45 VSS VDD 3 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=980 $Y=1010 $D=26
M46 3 VDD VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=1410 $Y=-840 $D=26
M47 3 VDD VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=1410 $Y=1010 $D=26
M48 VSS S[0] 5 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=3750 $Y=-840 $D=26
M49 VSS S[0] 5 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=3750 $Y=1010 $D=26
M50 5 S[0] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=4180 $Y=-840 $D=26
M51 5 S[0] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=4180 $Y=1010 $D=26
M52 VSS S[1] 7 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=6260 $Y=-840 $D=26
M53 VSS S[1] 7 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=6260 $Y=1010 $D=26
M54 7 S[1] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=6690 $Y=-840 $D=26
M55 7 S[1] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=6690 $Y=1010 $D=26
M56 VSS S[2] 9 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=9030 $Y=-840 $D=26
M57 VSS S[2] 9 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=9030 $Y=1010 $D=26
M58 9 S[2] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=9460 $Y=-840 $D=26
M59 9 S[2] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=9460 $Y=1010 $D=26
M60 VSS S[2] 9 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=11555 $Y=-840 $D=26
M61 VSS S[2] 9 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=11555 $Y=1010 $D=26
M62 9 S[2] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=11985 $Y=-840 $D=26
M63 9 S[2] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=11985 $Y=1010 $D=26
M64 VSS S[3] 11 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=14325 $Y=-840 $D=26
M65 VSS S[3] 11 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=14325 $Y=1010 $D=26
M66 11 S[3] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=14755 $Y=-840 $D=26
M67 11 S[3] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=14755 $Y=1010 $D=26
M68 VSS S[3] 11 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=16835 $Y=-840 $D=26
M69 VSS S[3] 11 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=16835 $Y=1010 $D=26
M70 11 S[3] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=17265 $Y=-840 $D=26
M71 11 S[3] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=17265 $Y=1010 $D=26
M72 VSS S[4] 13 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=19605 $Y=-840 $D=26
M73 VSS S[4] 13 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=19605 $Y=1010 $D=26
M74 13 S[4] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=20035 $Y=-840 $D=26
M75 13 S[4] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=20035 $Y=1010 $D=26
M76 VSS S[4] 13 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=22200 $Y=-840 $D=26
M77 VSS S[4] 13 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=22200 $Y=1010 $D=26
M78 13 S[4] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=22630 $Y=-840 $D=26
M79 13 S[4] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=22630 $Y=1010 $D=26
M80 VSS S[5] 16 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=24970 $Y=-840 $D=26
M81 VSS S[5] 16 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=24970 $Y=1010 $D=26
M82 16 S[5] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=25400 $Y=-840 $D=26
M83 16 S[5] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=25400 $Y=1010 $D=26
M84 VSS S[5] 16 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=27480 $Y=-840 $D=26
M85 VSS S[5] 16 VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=27480 $Y=1010 $D=26
M86 16 S[5] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=27910 $Y=-840 $D=26
M87 16 S[5] VSS VSS RFNPDHVT L=7E-08 W=4.6E-07 $X=27910 $Y=1010 $D=26
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PXA                                                                  *
*******************************************************************************
.SUBCKT qspi_data_info_32_memPXA VDD VSS PX[3] PX[2] PX[1] PX[0] A[0] A[1] CLK CLKX RDE


M0 29 19 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=115 $Y=3520 $D=0
M1 PX[0] 4 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=115 $Y=10345 $D=0
M2 9 CLKX 4 VSS N12LL L=6E-08 W=8.35E-07 $X=265 $Y=7855 $D=0
M3 VSS PX[0] 4 VSS N12LL L=6E-07 W=1.2E-07 $X=365 $Y=9535 $D=0
M4 19 12 VSS VSS N12LL L=6E-08 W=7E-07 $X=395 $Y=1550 $D=0
M5 9 5 29 VSS N12LL L=6E-08 W=7.5E-07 $X=405 $Y=3520 $D=0
M6 VSS 4 PX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=405 $Y=10345 $D=0
M7 4 CLKX 9 VSS N12LL L=6E-08 W=8.35E-07 $X=545 $Y=7855 $D=0
M8 VSS RDE 19 VSS N12LL L=6E-08 W=7E-07 $X=685 $Y=1550 $D=0
M9 30 5 9 VSS N12LL L=6E-08 W=7.5E-07 $X=695 $Y=3520 $D=0
M10 PX[0] 4 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=695 $Y=10345 $D=0
M11 9 CLKX 4 VSS N12LL L=6E-08 W=8.35E-07 $X=825 $Y=7855 $D=0
M12 10 RDE VSS VSS N12LL L=6E-08 W=5E-07 $X=975 $Y=1665 $D=0
M13 VSS 19 30 VSS N12LL L=6E-08 W=7.5E-07 $X=985 $Y=3520 $D=0
M14 VSS 4 PX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=985 $Y=10345 $D=0
M15 VSS 16 10 VSS N12LL L=6E-08 W=5E-07 $X=1265 $Y=1665 $D=0
M16 31 10 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1275 $Y=3520 $D=0
M17 PX[1] 13 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1275 $Y=10345 $D=0
M18 13 PX[1] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=1355 $Y=9535 $D=0
M19 13 CLKX 14 VSS N12LL L=6E-08 W=8.35E-07 $X=1435 $Y=7855 $D=0
M20 14 5 31 VSS N12LL L=6E-08 W=7.5E-07 $X=1565 $Y=3520 $D=0
M21 VSS 13 PX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1565 $Y=10345 $D=0
M22 14 CLKX 13 VSS N12LL L=6E-08 W=8.35E-07 $X=1715 $Y=7855 $D=0
M23 32 5 14 VSS N12LL L=6E-08 W=7.5E-07 $X=1855 $Y=3520 $D=0
M24 PX[1] 13 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1855 $Y=10345 $D=0
M25 VSS 16 12 VSS N12LL L=6E-08 W=4E-07 $X=1885 $Y=1550 $D=0
M26 13 CLKX 14 VSS N12LL L=6E-08 W=8.35E-07 $X=1995 $Y=7855 $D=0
M27 VSS 10 32 VSS N12LL L=6E-08 W=7.5E-07 $X=2145 $Y=3520 $D=0
M28 VSS 13 PX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=2145 $Y=10345 $D=0
M29 16 A[0] VSS VSS N12LL L=6E-08 W=4E-07 $X=2165 $Y=1550 $D=0
M30 33 10 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=2435 $Y=3520 $D=0
M31 PX[3] 17 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=2435 $Y=10345 $D=0
M32 21 CLKX 17 VSS N12LL L=6E-08 W=8.35E-07 $X=2585 $Y=7855 $D=0
M33 VSS PX[3] 17 VSS N12LL L=6E-07 W=1.2E-07 $X=2685 $Y=9535 $D=0
M34 21 18 33 VSS N12LL L=6E-08 W=7.5E-07 $X=2725 $Y=3520 $D=0
M35 VSS 17 PX[3] VSS N12LL L=6E-08 W=7.5E-07 $X=2725 $Y=10345 $D=0
M36 35 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=2795 $Y=1550 $D=0
M37 17 CLKX 21 VSS N12LL L=6E-08 W=8.35E-07 $X=2865 $Y=7855 $D=0
M38 34 18 21 VSS N12LL L=6E-08 W=7.5E-07 $X=3015 $Y=3520 $D=0
M39 PX[3] 17 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=3015 $Y=10345 $D=0
M40 21 CLKX 17 VSS N12LL L=6E-08 W=8.35E-07 $X=3145 $Y=7855 $D=0
M41 23 A[1] 35 VSS N12LL L=6E-08 W=4E-07 $X=3265 $Y=1550 $D=0
M42 VSS 10 34 VSS N12LL L=6E-08 W=7.5E-07 $X=3305 $Y=3520 $D=0
M43 VSS 17 PX[3] VSS N12LL L=6E-08 W=7.5E-07 $X=3305 $Y=10345 $D=0
M44 36 19 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=3595 $Y=3520 $D=0
M45 PX[2] 25 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=3595 $Y=10345 $D=0
M46 25 PX[2] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=3675 $Y=9535 $D=0
M47 25 CLKX 26 VSS N12LL L=6E-08 W=8.35E-07 $X=3755 $Y=7855 $D=0
M48 26 18 36 VSS N12LL L=6E-08 W=7.5E-07 $X=3885 $Y=3520 $D=0
M49 VSS 25 PX[2] VSS N12LL L=6E-08 W=7.5E-07 $X=3885 $Y=10345 $D=0
M50 VSS 23 18 VSS N12LL L=6E-08 W=7E-07 $X=3895 $Y=1550 $D=0
M51 26 CLKX 25 VSS N12LL L=6E-08 W=8.35E-07 $X=4035 $Y=7855 $D=0
M52 37 18 26 VSS N12LL L=6E-08 W=7.5E-07 $X=4175 $Y=3520 $D=0
M53 PX[2] 25 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=4175 $Y=10345 $D=0
M54 5 18 VSS VSS N12LL L=6E-08 W=7E-07 $X=4185 $Y=1550 $D=0
M55 25 CLKX 26 VSS N12LL L=6E-08 W=8.35E-07 $X=4315 $Y=7855 $D=0
M56 VSS 19 37 VSS N12LL L=6E-08 W=7.5E-07 $X=4465 $Y=3520 $D=0
M57 VSS 25 PX[2] VSS N12LL L=6E-08 W=7.5E-07 $X=4465 $Y=10345 $D=0
M58 9 19 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=115 $Y=4770 $D=1
M59 PX[0] 4 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=115 $Y=11695 $D=1
M60 9 CLK 4 VDD P12LL L=6E-08 W=8.3E-07 $X=265 $Y=6525 $D=1
M61 38 12 19 VDD P12LL L=6E-08 W=1.4E-06 $X=395 $Y=-450 $D=1
M62 VDD 5 9 VDD P12LL L=6E-08 W=7.5E-07 $X=405 $Y=4770 $D=1
M63 VDD 4 PX[0] VDD P12LL L=6E-08 W=1.75E-06 $X=405 $Y=11695 $D=1
M64 4 CLK 9 VDD P12LL L=6E-08 W=8.3E-07 $X=545 $Y=6525 $D=1
M65 VDD PX[0] 4 VDD P12LL L=3E-07 W=1.2E-07 $X=615 $Y=14130 $D=1
M66 VDD RDE 38 VDD P12LL L=6E-08 W=1.4E-06 $X=685 $Y=-450 $D=1
M67 9 5 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=695 $Y=4770 $D=1
M68 PX[0] 4 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=695 $Y=11695 $D=1
M69 9 CLK 4 VDD P12LL L=6E-08 W=8.3E-07 $X=825 $Y=6525 $D=1
M70 39 RDE VDD VDD P12LL L=6E-08 W=7E-07 $X=975 $Y=250 $D=1
M71 VDD 19 9 VDD P12LL L=6E-08 W=7.5E-07 $X=985 $Y=4770 $D=1
M72 VDD 4 PX[0] VDD P12LL L=6E-08 W=1.75E-06 $X=985 $Y=11695 $D=1
M73 10 16 39 VDD P12LL L=6E-08 W=7E-07 $X=1265 $Y=250 $D=1
M74 14 10 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=1275 $Y=4770 $D=1
M75 PX[1] 13 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=1275 $Y=11695 $D=1
M76 13 PX[1] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=1405 $Y=14130 $D=1
M77 13 CLK 14 VDD P12LL L=6E-08 W=8.3E-07 $X=1435 $Y=6525 $D=1
M78 VDD 5 14 VDD P12LL L=6E-08 W=7.5E-07 $X=1565 $Y=4770 $D=1
M79 VDD 13 PX[1] VDD P12LL L=6E-08 W=1.75E-06 $X=1565 $Y=11695 $D=1
M80 14 CLK 13 VDD P12LL L=6E-08 W=8.3E-07 $X=1715 $Y=6525 $D=1
M81 14 5 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=1855 $Y=4770 $D=1
M82 PX[1] 13 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=1855 $Y=11695 $D=1
M83 VDD 16 12 VDD P12LL L=6E-08 W=4E-07 $X=1885 $Y=400 $D=1
M84 13 CLK 14 VDD P12LL L=6E-08 W=8.3E-07 $X=1995 $Y=6525 $D=1
M85 VDD 10 14 VDD P12LL L=6E-08 W=7.5E-07 $X=2145 $Y=4770 $D=1
M86 VDD 13 PX[1] VDD P12LL L=6E-08 W=1.75E-06 $X=2145 $Y=11695 $D=1
M87 16 A[0] VDD VDD P12LL L=6E-08 W=4E-07 $X=2165 $Y=400 $D=1
M88 21 10 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=2435 $Y=4770 $D=1
M89 PX[3] 17 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=2435 $Y=11695 $D=1
M90 21 CLK 17 VDD P12LL L=6E-08 W=8.3E-07 $X=2585 $Y=6525 $D=1
M91 VDD 18 21 VDD P12LL L=6E-08 W=7.5E-07 $X=2725 $Y=4770 $D=1
M92 VDD 17 PX[3] VDD P12LL L=6E-08 W=1.75E-06 $X=2725 $Y=11695 $D=1
M93 17 CLK 21 VDD P12LL L=6E-08 W=8.3E-07 $X=2865 $Y=6525 $D=1
M94 VDD PX[3] 17 VDD P12LL L=3E-07 W=1.2E-07 $X=2935 $Y=14130 $D=1
M95 41 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=2995 $Y=485 $D=1
M96 21 18 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=3015 $Y=4770 $D=1
M97 PX[3] 17 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=3015 $Y=11695 $D=1
M98 21 CLK 17 VDD P12LL L=6E-08 W=8.3E-07 $X=3145 $Y=6525 $D=1
M99 23 A[1] 41 VDD P12LL L=6E-08 W=4E-07 $X=3265 $Y=485 $D=1
M100 VDD 10 21 VDD P12LL L=6E-08 W=7.5E-07 $X=3305 $Y=4770 $D=1
M101 VDD 17 PX[3] VDD P12LL L=6E-08 W=1.75E-06 $X=3305 $Y=11695 $D=1
M102 26 19 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=3595 $Y=4770 $D=1
M103 PX[2] 25 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=3595 $Y=11695 $D=1
M104 25 PX[2] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=3725 $Y=14130 $D=1
M105 25 CLK 26 VDD P12LL L=6E-08 W=8.3E-07 $X=3755 $Y=6525 $D=1
M106 VDD 18 26 VDD P12LL L=6E-08 W=7.5E-07 $X=3885 $Y=4770 $D=1
M107 VDD 25 PX[2] VDD P12LL L=6E-08 W=1.75E-06 $X=3885 $Y=11695 $D=1
M108 VDD 23 18 VDD P12LL L=6E-08 W=1.4E-06 $X=3895 $Y=-450 $D=1
M109 26 CLK 25 VDD P12LL L=6E-08 W=8.3E-07 $X=4035 $Y=6525 $D=1
M110 26 18 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=4175 $Y=4770 $D=1
M111 PX[2] 25 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=4175 $Y=11695 $D=1
M112 5 18 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=4185 $Y=-450 $D=1
M113 25 CLK 26 VDD P12LL L=6E-08 W=8.3E-07 $X=4315 $Y=6525 $D=1
M114 VDD 19 26 VDD P12LL L=6E-08 W=7.5E-07 $X=4465 $Y=4770 $D=1
M115 VDD 25 PX[2] VDD P12LL L=6E-08 W=1.75E-06 $X=4465 $Y=11695 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: FPREDEC                                                              *
*******************************************************************************
.SUBCKT qspi_data_info_32_memFPREDEC VDD VSS FCKX[7] FCKX[6] FCKX[5] FCKX[4] FCKX[3] FCKX[2] FCKX[1] FCKX[0]
+A[0] A[1] A[2] CLK CLKX WLCKX


M0 6 4 VSS VSS N12LL L=6E-08 W=4E-07 $X=115 $Y=10310 $D=0
M1 FCKX[3] 6 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=115 $Y=14130 $D=0
M2 23 45 VSS VSS N12LL L=6E-08 W=5E-07 $X=255 $Y=140 $D=0
M3 7 CLKX 4 VSS N12LL L=6E-08 W=5E-07 $X=275 $Y=6170 $D=0
M4 VSS 6 4 VSS N12LL L=6E-07 W=1.2E-07 $X=365 $Y=11505 $D=0
M5 VSS 4 6 VSS N12LL L=6E-08 W=4E-07 $X=405 $Y=10310 $D=0
M6 WLCKX 6 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=405 $Y=14130 $D=0
M7 57 5 7 VSS N12LL L=6E-08 W=1E-06 $X=505 $Y=4625 $D=0
M8 VSS 45 23 VSS N12LL L=6E-08 W=5E-07 $X=545 $Y=140 $D=0
M9 4 CLKX 7 VSS N12LL L=6E-08 W=5E-07 $X=545 $Y=6170 $D=0
M10 6 4 VSS VSS N12LL L=6E-08 W=4E-07 $X=695 $Y=10310 $D=0
M11 FCKX[3] 6 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=695 $Y=14130 $D=0
M12 58 10 57 VSS N12LL L=6E-08 W=1E-06 $X=745 $Y=4625 $D=0
M13 7 CLKX 4 VSS N12LL L=6E-08 W=5E-07 $X=825 $Y=6170 $D=0
M14 45 11 VSS VSS N12LL L=6E-08 W=5E-07 $X=835 $Y=140 $D=0
M15 VSS 23 58 VSS N12LL L=6E-08 W=1E-06 $X=985 $Y=4625 $D=0
M16 VSS 4 6 VSS N12LL L=6E-08 W=4E-07 $X=985 $Y=10310 $D=0
M17 WLCKX 6 FCKX[3] VSS N12LL L=6E-08 W=1.25E-06 $X=985 $Y=14130 $D=0
M18 VSS 11 45 VSS N12LL L=6E-08 W=5E-07 $X=1125 $Y=140 $D=0
M19 59 23 VSS VSS N12LL L=6E-08 W=1E-06 $X=1275 $Y=4625 $D=0
M20 12 14 VSS VSS N12LL L=6E-08 W=4E-07 $X=1275 $Y=10310 $D=0
M21 FCKX[2] 12 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=1275 $Y=14130 $D=0
M22 14 12 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=1355 $Y=11505 $D=0
M23 14 CLKX 13 VSS N12LL L=6E-08 W=5E-07 $X=1435 $Y=6170 $D=0
M24 60 10 59 VSS N12LL L=6E-08 W=1E-06 $X=1515 $Y=4625 $D=0
M25 VSS 14 12 VSS N12LL L=6E-08 W=4E-07 $X=1565 $Y=10310 $D=0
M26 WLCKX 12 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=1565 $Y=14130 $D=0
M27 13 CLKX 14 VSS N12LL L=6E-08 W=5E-07 $X=1715 $Y=6170 $D=0
M28 61 A[2] 11 VSS N12LL L=6E-08 W=4E-07 $X=1755 $Y=160 $D=0
M29 13 18 60 VSS N12LL L=6E-08 W=1E-06 $X=1755 $Y=4625 $D=0
M30 12 14 VSS VSS N12LL L=6E-08 W=4E-07 $X=1855 $Y=10310 $D=0
M31 FCKX[2] 12 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=1855 $Y=14130 $D=0
M32 14 CLKX 13 VSS N12LL L=6E-08 W=5E-07 $X=1985 $Y=6170 $D=0
M33 VSS VDD 61 VSS N12LL L=3E-07 W=4E-07 $X=2015 $Y=160 $D=0
M34 VSS 14 12 VSS N12LL L=6E-08 W=4E-07 $X=2145 $Y=10310 $D=0
M35 WLCKX 12 FCKX[2] VSS N12LL L=6E-08 W=1.25E-06 $X=2145 $Y=14130 $D=0
M36 21 19 VSS VSS N12LL L=6E-08 W=4E-07 $X=2435 $Y=10310 $D=0
M37 FCKX[0] 21 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=2435 $Y=14130 $D=0
M38 22 CLKX 19 VSS N12LL L=6E-08 W=5E-07 $X=2595 $Y=6170 $D=0
M39 VSS 21 19 VSS N12LL L=6E-07 W=1.2E-07 $X=2685 $Y=11505 $D=0
M40 VSS 19 21 VSS N12LL L=6E-08 W=4E-07 $X=2725 $Y=10310 $D=0
M41 WLCKX 21 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=2725 $Y=14130 $D=0
M42 62 18 22 VSS N12LL L=6E-08 W=1E-06 $X=2825 $Y=4625 $D=0
M43 19 CLKX 22 VSS N12LL L=6E-08 W=5E-07 $X=2865 $Y=6170 $D=0
M44 21 19 VSS VSS N12LL L=6E-08 W=4E-07 $X=3015 $Y=10310 $D=0
M45 FCKX[0] 21 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=3015 $Y=14130 $D=0
M46 63 53 62 VSS N12LL L=6E-08 W=1E-06 $X=3065 $Y=4625 $D=0
M47 22 CLKX 19 VSS N12LL L=6E-08 W=5E-07 $X=3145 $Y=6170 $D=0
M48 VSS 23 63 VSS N12LL L=6E-08 W=1E-06 $X=3305 $Y=4625 $D=0
M49 VSS 19 21 VSS N12LL L=6E-08 W=4E-07 $X=3305 $Y=10310 $D=0
M50 WLCKX 21 FCKX[0] VSS N12LL L=6E-08 W=1.25E-06 $X=3305 $Y=14130 $D=0
M51 64 23 VSS VSS N12LL L=6E-08 W=1E-06 $X=3595 $Y=4625 $D=0
M52 26 27 VSS VSS N12LL L=6E-08 W=4E-07 $X=3595 $Y=10310 $D=0
M53 FCKX[1] 26 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=3595 $Y=14130 $D=0
M54 27 26 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=3675 $Y=11505 $D=0
M55 27 CLKX 28 VSS N12LL L=6E-08 W=5E-07 $X=3755 $Y=6170 $D=0
M56 65 53 64 VSS N12LL L=6E-08 W=1E-06 $X=3835 $Y=4625 $D=0
M57 VSS 27 26 VSS N12LL L=6E-08 W=4E-07 $X=3885 $Y=10310 $D=0
M58 WLCKX 26 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=3885 $Y=14130 $D=0
M59 28 CLKX 27 VSS N12LL L=6E-08 W=5E-07 $X=4035 $Y=6170 $D=0
M60 66 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=4065 $Y=160 $D=0
M61 28 5 65 VSS N12LL L=6E-08 W=1E-06 $X=4075 $Y=4625 $D=0
M62 26 27 VSS VSS N12LL L=6E-08 W=4E-07 $X=4175 $Y=10310 $D=0
M63 FCKX[1] 26 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=4175 $Y=14130 $D=0
M64 27 CLKX 28 VSS N12LL L=6E-08 W=5E-07 $X=4305 $Y=6170 $D=0
M65 VSS 27 26 VSS N12LL L=6E-08 W=4E-07 $X=4465 $Y=10310 $D=0
M66 WLCKX 26 FCKX[1] VSS N12LL L=6E-08 W=1.25E-06 $X=4465 $Y=14130 $D=0
M67 32 A[0] 66 VSS N12LL L=6E-08 W=4E-07 $X=4565 $Y=160 $D=0
M68 33 31 VSS VSS N12LL L=6E-08 W=4E-07 $X=4755 $Y=10310 $D=0
M69 FCKX[7] 33 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=4755 $Y=14130 $D=0
M70 34 CLKX 31 VSS N12LL L=6E-08 W=5E-07 $X=4915 $Y=6170 $D=0
M71 VSS 33 31 VSS N12LL L=6E-07 W=1.2E-07 $X=5005 $Y=11505 $D=0
M72 VSS 31 33 VSS N12LL L=6E-08 W=4E-07 $X=5045 $Y=10310 $D=0
M73 WLCKX 33 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=5045 $Y=14130 $D=0
M74 67 5 34 VSS N12LL L=6E-08 W=1E-06 $X=5145 $Y=4625 $D=0
M75 31 CLKX 34 VSS N12LL L=6E-08 W=5E-07 $X=5185 $Y=6170 $D=0
M76 5 32 VSS VSS N12LL L=6E-08 W=5E-07 $X=5195 $Y=140 $D=0
M77 33 31 VSS VSS N12LL L=6E-08 W=4E-07 $X=5335 $Y=10310 $D=0
M78 FCKX[7] 33 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=5335 $Y=14130 $D=0
M79 68 10 67 VSS N12LL L=6E-08 W=1E-06 $X=5385 $Y=4625 $D=0
M80 34 CLKX 31 VSS N12LL L=6E-08 W=5E-07 $X=5465 $Y=6170 $D=0
M81 VSS 32 5 VSS N12LL L=6E-08 W=5E-07 $X=5485 $Y=140 $D=0
M82 VSS 45 68 VSS N12LL L=6E-08 W=1E-06 $X=5625 $Y=4625 $D=0
M83 VSS 31 33 VSS N12LL L=6E-08 W=4E-07 $X=5625 $Y=10310 $D=0
M84 WLCKX 33 FCKX[7] VSS N12LL L=6E-08 W=1.25E-06 $X=5625 $Y=14130 $D=0
M85 18 5 VSS VSS N12LL L=6E-08 W=5E-07 $X=5775 $Y=140 $D=0
M86 69 45 VSS VSS N12LL L=6E-08 W=1E-06 $X=5915 $Y=4625 $D=0
M87 36 38 VSS VSS N12LL L=6E-08 W=4E-07 $X=5915 $Y=10310 $D=0
M88 FCKX[6] 36 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=5915 $Y=14130 $D=0
M89 38 36 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=5995 $Y=11505 $D=0
M90 VSS 5 18 VSS N12LL L=6E-08 W=5E-07 $X=6065 $Y=140 $D=0
M91 38 CLKX 37 VSS N12LL L=6E-08 W=5E-07 $X=6075 $Y=6170 $D=0
M92 70 10 69 VSS N12LL L=6E-08 W=1E-06 $X=6155 $Y=4625 $D=0
M93 VSS 38 36 VSS N12LL L=6E-08 W=4E-07 $X=6205 $Y=10310 $D=0
M94 WLCKX 36 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=6205 $Y=14130 $D=0
M95 37 CLKX 38 VSS N12LL L=6E-08 W=5E-07 $X=6355 $Y=6170 $D=0
M96 37 18 70 VSS N12LL L=6E-08 W=1E-06 $X=6395 $Y=4625 $D=0
M97 36 38 VSS VSS N12LL L=6E-08 W=4E-07 $X=6495 $Y=10310 $D=0
M98 FCKX[6] 36 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=6495 $Y=14130 $D=0
M99 38 CLKX 37 VSS N12LL L=6E-08 W=5E-07 $X=6625 $Y=6170 $D=0
M100 VSS 38 36 VSS N12LL L=6E-08 W=4E-07 $X=6785 $Y=10310 $D=0
M101 WLCKX 36 FCKX[6] VSS N12LL L=6E-08 W=1.25E-06 $X=6785 $Y=14130 $D=0
M102 43 42 VSS VSS N12LL L=6E-08 W=4E-07 $X=7075 $Y=10310 $D=0
M103 FCKX[4] 43 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=7075 $Y=14130 $D=0
M104 71 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=7105 $Y=160 $D=0
M105 44 CLKX 42 VSS N12LL L=6E-08 W=5E-07 $X=7235 $Y=6170 $D=0
M106 VSS 43 42 VSS N12LL L=6E-07 W=1.2E-07 $X=7325 $Y=11505 $D=0
M107 VSS 42 43 VSS N12LL L=6E-08 W=4E-07 $X=7365 $Y=10310 $D=0
M108 WLCKX 43 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=7365 $Y=14130 $D=0
M109 72 18 44 VSS N12LL L=6E-08 W=1E-06 $X=7465 $Y=4625 $D=0
M110 42 CLKX 44 VSS N12LL L=6E-08 W=5E-07 $X=7505 $Y=6170 $D=0
M111 47 A[1] 71 VSS N12LL L=6E-08 W=4E-07 $X=7605 $Y=160 $D=0
M112 43 42 VSS VSS N12LL L=6E-08 W=4E-07 $X=7655 $Y=10310 $D=0
M113 FCKX[4] 43 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=7655 $Y=14130 $D=0
M114 73 53 72 VSS N12LL L=6E-08 W=1E-06 $X=7705 $Y=4625 $D=0
M115 44 CLKX 42 VSS N12LL L=6E-08 W=5E-07 $X=7785 $Y=6170 $D=0
M116 VSS 45 73 VSS N12LL L=6E-08 W=1E-06 $X=7945 $Y=4625 $D=0
M117 VSS 42 43 VSS N12LL L=6E-08 W=4E-07 $X=7945 $Y=10310 $D=0
M118 WLCKX 43 FCKX[4] VSS N12LL L=6E-08 W=1.25E-06 $X=7945 $Y=14130 $D=0
M119 10 47 VSS VSS N12LL L=6E-08 W=5E-07 $X=8235 $Y=140 $D=0
M120 74 45 VSS VSS N12LL L=6E-08 W=1E-06 $X=8235 $Y=4625 $D=0
M121 48 49 VSS VSS N12LL L=6E-08 W=4E-07 $X=8235 $Y=10310 $D=0
M122 FCKX[5] 48 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=8235 $Y=14130 $D=0
M123 49 48 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=8315 $Y=11505 $D=0
M124 49 CLKX 50 VSS N12LL L=6E-08 W=5E-07 $X=8395 $Y=6170 $D=0
M125 75 53 74 VSS N12LL L=6E-08 W=1E-06 $X=8475 $Y=4625 $D=0
M126 VSS 47 10 VSS N12LL L=6E-08 W=5E-07 $X=8525 $Y=140 $D=0
M127 VSS 49 48 VSS N12LL L=6E-08 W=4E-07 $X=8525 $Y=10310 $D=0
M128 WLCKX 48 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=8525 $Y=14130 $D=0
M129 50 CLKX 49 VSS N12LL L=6E-08 W=5E-07 $X=8675 $Y=6170 $D=0
M130 50 5 75 VSS N12LL L=6E-08 W=1E-06 $X=8715 $Y=4625 $D=0
M131 53 10 VSS VSS N12LL L=6E-08 W=5E-07 $X=8815 $Y=140 $D=0
M132 48 49 VSS VSS N12LL L=6E-08 W=4E-07 $X=8815 $Y=10310 $D=0
M133 FCKX[5] 48 WLCKX VSS N12LL L=6E-08 W=1.25E-06 $X=8815 $Y=14130 $D=0
M134 49 CLKX 50 VSS N12LL L=6E-08 W=5E-07 $X=8945 $Y=6170 $D=0
M135 VSS 10 53 VSS N12LL L=6E-08 W=5E-07 $X=9105 $Y=140 $D=0
M136 VSS 49 48 VSS N12LL L=6E-08 W=4E-07 $X=9105 $Y=10310 $D=0
M137 WLCKX 48 FCKX[5] VSS N12LL L=6E-08 W=1.25E-06 $X=9105 $Y=14130 $D=0
M138 6 4 VDD VDD P12LL L=6E-08 W=4E-07 $X=115 $Y=9125 $D=1
M139 FCKX[3] 4 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=115 $Y=12320 $D=1
M140 FCKX[3] 6 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=115 $Y=15880 $D=1
M141 23 45 VDD VDD P12LL L=6E-08 W=1E-06 $X=255 $Y=1195 $D=1
M142 7 CLK 4 VDD P12LL L=6E-08 W=5E-07 $X=275 $Y=7170 $D=1
M143 VDD 5 7 VDD P12LL L=6E-08 W=1E-06 $X=405 $Y=3025 $D=1
M144 VDD 4 6 VDD P12LL L=6E-08 W=4E-07 $X=405 $Y=9125 $D=1
M145 WLCKX 4 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=405 $Y=12320 $D=1
M146 VDD 6 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=405 $Y=15880 $D=1
M147 VDD 45 23 VDD P12LL L=6E-08 W=1E-06 $X=545 $Y=1195 $D=1
M148 4 CLK 7 VDD P12LL L=6E-08 W=5E-07 $X=545 $Y=7170 $D=1
M149 VDD 6 4 VDD P12LL L=3E-07 W=1.2E-07 $X=655 $Y=8285 $D=1
M150 7 10 VDD VDD P12LL L=6E-08 W=1E-06 $X=695 $Y=3025 $D=1
M151 6 4 VDD VDD P12LL L=6E-08 W=4E-07 $X=695 $Y=9125 $D=1
M152 FCKX[3] 4 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=695 $Y=12320 $D=1
M153 FCKX[3] 6 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=695 $Y=15880 $D=1
M154 7 CLK 4 VDD P12LL L=6E-08 W=5E-07 $X=825 $Y=7170 $D=1
M155 45 11 VDD VDD P12LL L=6E-08 W=1E-06 $X=835 $Y=1195 $D=1
M156 VDD 23 7 VDD P12LL L=6E-08 W=1E-06 $X=985 $Y=3025 $D=1
M157 VDD 4 6 VDD P12LL L=6E-08 W=4E-07 $X=985 $Y=9125 $D=1
M158 WLCKX 4 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=985 $Y=12320 $D=1
M159 VDD 6 FCKX[3] VDD P12LL L=6E-08 W=1.25E-06 $X=985 $Y=15880 $D=1
M160 VDD 11 45 VDD P12LL L=6E-08 W=1E-06 $X=1125 $Y=1195 $D=1
M161 13 23 VDD VDD P12LL L=6E-08 W=1E-06 $X=1275 $Y=3025 $D=1
M162 12 14 VDD VDD P12LL L=6E-08 W=4E-07 $X=1275 $Y=9125 $D=1
M163 FCKX[2] 14 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=1275 $Y=12320 $D=1
M164 FCKX[2] 12 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=1275 $Y=15880 $D=1
M165 14 12 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=1365 $Y=8285 $D=1
M166 14 CLK 13 VDD P12LL L=6E-08 W=5E-07 $X=1435 $Y=7170 $D=1
M167 VDD 10 13 VDD P12LL L=6E-08 W=1E-06 $X=1565 $Y=3025 $D=1
M168 VDD 14 12 VDD P12LL L=6E-08 W=4E-07 $X=1565 $Y=9125 $D=1
M169 WLCKX 14 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=1565 $Y=12320 $D=1
M170 VDD 12 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=1565 $Y=15880 $D=1
M171 13 CLK 14 VDD P12LL L=6E-08 W=5E-07 $X=1715 $Y=7170 $D=1
M172 77 A[2] 11 VDD P12LL L=6E-08 W=4E-07 $X=1755 $Y=1245 $D=1
M173 13 18 VDD VDD P12LL L=6E-08 W=1E-06 $X=1855 $Y=3025 $D=1
M174 12 14 VDD VDD P12LL L=6E-08 W=4E-07 $X=1855 $Y=9125 $D=1
M175 FCKX[2] 14 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=1855 $Y=12320 $D=1
M176 FCKX[2] 12 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=1855 $Y=15880 $D=1
M177 VDD VSS 77 VDD P12LL L=1E-07 W=4E-07 $X=1985 $Y=1245 $D=1
M178 14 CLK 13 VDD P12LL L=6E-08 W=5E-07 $X=1985 $Y=7170 $D=1
M179 VDD 14 12 VDD P12LL L=6E-08 W=4E-07 $X=2145 $Y=9125 $D=1
M180 WLCKX 14 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=2145 $Y=12320 $D=1
M181 VDD 12 FCKX[2] VDD P12LL L=6E-08 W=1.25E-06 $X=2145 $Y=15880 $D=1
M182 21 19 VDD VDD P12LL L=6E-08 W=4E-07 $X=2435 $Y=9125 $D=1
M183 FCKX[0] 19 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=2435 $Y=12320 $D=1
M184 FCKX[0] 21 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=2435 $Y=15880 $D=1
M185 22 CLK 19 VDD P12LL L=6E-08 W=5E-07 $X=2595 $Y=7170 $D=1
M186 VDD 18 22 VDD P12LL L=6E-08 W=1E-06 $X=2725 $Y=3025 $D=1
M187 VDD 19 21 VDD P12LL L=6E-08 W=4E-07 $X=2725 $Y=9125 $D=1
M188 WLCKX 19 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=2725 $Y=12320 $D=1
M189 VDD 21 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=2725 $Y=15880 $D=1
M190 19 CLK 22 VDD P12LL L=6E-08 W=5E-07 $X=2865 $Y=7170 $D=1
M191 VDD 21 19 VDD P12LL L=3E-07 W=1.2E-07 $X=2975 $Y=8285 $D=1
M192 22 53 VDD VDD P12LL L=6E-08 W=1E-06 $X=3015 $Y=3025 $D=1
M193 21 19 VDD VDD P12LL L=6E-08 W=4E-07 $X=3015 $Y=9125 $D=1
M194 FCKX[0] 19 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=3015 $Y=12320 $D=1
M195 FCKX[0] 21 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=3015 $Y=15880 $D=1
M196 22 CLK 19 VDD P12LL L=6E-08 W=5E-07 $X=3145 $Y=7170 $D=1
M197 VDD 23 22 VDD P12LL L=6E-08 W=1E-06 $X=3305 $Y=3025 $D=1
M198 VDD 19 21 VDD P12LL L=6E-08 W=4E-07 $X=3305 $Y=9125 $D=1
M199 WLCKX 19 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=3305 $Y=12320 $D=1
M200 VDD 21 FCKX[0] VDD P12LL L=6E-08 W=1.25E-06 $X=3305 $Y=15880 $D=1
M201 28 23 VDD VDD P12LL L=6E-08 W=1E-06 $X=3595 $Y=3025 $D=1
M202 26 27 VDD VDD P12LL L=6E-08 W=4E-07 $X=3595 $Y=9125 $D=1
M203 FCKX[1] 27 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=3595 $Y=12320 $D=1
M204 FCKX[1] 26 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=3595 $Y=15880 $D=1
M205 27 26 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=3685 $Y=8285 $D=1
M206 27 CLK 28 VDD P12LL L=6E-08 W=5E-07 $X=3755 $Y=7170 $D=1
M207 VDD 53 28 VDD P12LL L=6E-08 W=1E-06 $X=3885 $Y=3025 $D=1
M208 VDD 27 26 VDD P12LL L=6E-08 W=4E-07 $X=3885 $Y=9125 $D=1
M209 WLCKX 27 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=3885 $Y=12320 $D=1
M210 VDD 26 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=3885 $Y=15880 $D=1
M211 28 CLK 27 VDD P12LL L=6E-08 W=5E-07 $X=4035 $Y=7170 $D=1
M212 28 5 VDD VDD P12LL L=6E-08 W=1E-06 $X=4175 $Y=3025 $D=1
M213 26 27 VDD VDD P12LL L=6E-08 W=4E-07 $X=4175 $Y=9125 $D=1
M214 FCKX[1] 27 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=4175 $Y=12320 $D=1
M215 FCKX[1] 26 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=4175 $Y=15880 $D=1
M216 78 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=4295 $Y=1245 $D=1
M217 27 CLK 28 VDD P12LL L=6E-08 W=5E-07 $X=4305 $Y=7170 $D=1
M218 VDD 27 26 VDD P12LL L=6E-08 W=4E-07 $X=4465 $Y=9125 $D=1
M219 WLCKX 27 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=4465 $Y=12320 $D=1
M220 VDD 26 FCKX[1] VDD P12LL L=6E-08 W=1.25E-06 $X=4465 $Y=15880 $D=1
M221 32 A[0] 78 VDD P12LL L=6E-08 W=4E-07 $X=4565 $Y=1245 $D=1
M222 33 31 VDD VDD P12LL L=6E-08 W=4E-07 $X=4755 $Y=9125 $D=1
M223 FCKX[7] 31 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=4755 $Y=12320 $D=1
M224 FCKX[7] 33 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=4755 $Y=15880 $D=1
M225 34 CLK 31 VDD P12LL L=6E-08 W=5E-07 $X=4915 $Y=7170 $D=1
M226 VDD 5 34 VDD P12LL L=6E-08 W=1E-06 $X=5045 $Y=3025 $D=1
M227 VDD 31 33 VDD P12LL L=6E-08 W=4E-07 $X=5045 $Y=9125 $D=1
M228 WLCKX 31 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=5045 $Y=12320 $D=1
M229 VDD 33 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=5045 $Y=15880 $D=1
M230 31 CLK 34 VDD P12LL L=6E-08 W=5E-07 $X=5185 $Y=7170 $D=1
M231 5 32 VDD VDD P12LL L=6E-08 W=1E-06 $X=5195 $Y=1195 $D=1
M232 VDD 33 31 VDD P12LL L=3E-07 W=1.2E-07 $X=5295 $Y=8285 $D=1
M233 34 10 VDD VDD P12LL L=6E-08 W=1E-06 $X=5335 $Y=3025 $D=1
M234 33 31 VDD VDD P12LL L=6E-08 W=4E-07 $X=5335 $Y=9125 $D=1
M235 FCKX[7] 31 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=5335 $Y=12320 $D=1
M236 FCKX[7] 33 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5335 $Y=15880 $D=1
M237 34 CLK 31 VDD P12LL L=6E-08 W=5E-07 $X=5465 $Y=7170 $D=1
M238 VDD 32 5 VDD P12LL L=6E-08 W=1E-06 $X=5485 $Y=1195 $D=1
M239 VDD 45 34 VDD P12LL L=6E-08 W=1E-06 $X=5625 $Y=3025 $D=1
M240 VDD 31 33 VDD P12LL L=6E-08 W=4E-07 $X=5625 $Y=9125 $D=1
M241 WLCKX 31 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=5625 $Y=12320 $D=1
M242 VDD 33 FCKX[7] VDD P12LL L=6E-08 W=1.25E-06 $X=5625 $Y=15880 $D=1
M243 18 5 VDD VDD P12LL L=6E-08 W=1E-06 $X=5775 $Y=1195 $D=1
M244 37 45 VDD VDD P12LL L=6E-08 W=1E-06 $X=5915 $Y=3025 $D=1
M245 36 38 VDD VDD P12LL L=6E-08 W=4E-07 $X=5915 $Y=9125 $D=1
M246 FCKX[6] 38 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=5915 $Y=12320 $D=1
M247 FCKX[6] 36 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5915 $Y=15880 $D=1
M248 38 36 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=6005 $Y=8285 $D=1
M249 VDD 5 18 VDD P12LL L=6E-08 W=1E-06 $X=6065 $Y=1195 $D=1
M250 38 CLK 37 VDD P12LL L=6E-08 W=5E-07 $X=6075 $Y=7170 $D=1
M251 VDD 10 37 VDD P12LL L=6E-08 W=1E-06 $X=6205 $Y=3025 $D=1
M252 VDD 38 36 VDD P12LL L=6E-08 W=4E-07 $X=6205 $Y=9125 $D=1
M253 WLCKX 38 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=6205 $Y=12320 $D=1
M254 VDD 36 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=6205 $Y=15880 $D=1
M255 37 CLK 38 VDD P12LL L=6E-08 W=5E-07 $X=6355 $Y=7170 $D=1
M256 37 18 VDD VDD P12LL L=6E-08 W=1E-06 $X=6495 $Y=3025 $D=1
M257 36 38 VDD VDD P12LL L=6E-08 W=4E-07 $X=6495 $Y=9125 $D=1
M258 FCKX[6] 38 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=6495 $Y=12320 $D=1
M259 FCKX[6] 36 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=6495 $Y=15880 $D=1
M260 38 CLK 37 VDD P12LL L=6E-08 W=5E-07 $X=6625 $Y=7170 $D=1
M261 VDD 38 36 VDD P12LL L=6E-08 W=4E-07 $X=6785 $Y=9125 $D=1
M262 WLCKX 38 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=6785 $Y=12320 $D=1
M263 VDD 36 FCKX[6] VDD P12LL L=6E-08 W=1.25E-06 $X=6785 $Y=15880 $D=1
M264 43 42 VDD VDD P12LL L=6E-08 W=4E-07 $X=7075 $Y=9125 $D=1
M265 FCKX[4] 42 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=7075 $Y=12320 $D=1
M266 FCKX[4] 43 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=7075 $Y=15880 $D=1
M267 44 CLK 42 VDD P12LL L=6E-08 W=5E-07 $X=7235 $Y=7170 $D=1
M268 79 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=7335 $Y=1245 $D=1
M269 VDD 18 44 VDD P12LL L=6E-08 W=1E-06 $X=7365 $Y=3025 $D=1
M270 VDD 42 43 VDD P12LL L=6E-08 W=4E-07 $X=7365 $Y=9125 $D=1
M271 WLCKX 42 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=7365 $Y=12320 $D=1
M272 VDD 43 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=7365 $Y=15880 $D=1
M273 42 CLK 44 VDD P12LL L=6E-08 W=5E-07 $X=7505 $Y=7170 $D=1
M274 47 A[1] 79 VDD P12LL L=6E-08 W=4E-07 $X=7605 $Y=1245 $D=1
M275 VDD 43 42 VDD P12LL L=3E-07 W=1.2E-07 $X=7615 $Y=8285 $D=1
M276 44 53 VDD VDD P12LL L=6E-08 W=1E-06 $X=7655 $Y=3025 $D=1
M277 43 42 VDD VDD P12LL L=6E-08 W=4E-07 $X=7655 $Y=9125 $D=1
M278 FCKX[4] 42 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=7655 $Y=12320 $D=1
M279 FCKX[4] 43 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=7655 $Y=15880 $D=1
M280 44 CLK 42 VDD P12LL L=6E-08 W=5E-07 $X=7785 $Y=7170 $D=1
M281 VDD 45 44 VDD P12LL L=6E-08 W=1E-06 $X=7945 $Y=3025 $D=1
M282 VDD 42 43 VDD P12LL L=6E-08 W=4E-07 $X=7945 $Y=9125 $D=1
M283 WLCKX 42 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=7945 $Y=12320 $D=1
M284 VDD 43 FCKX[4] VDD P12LL L=6E-08 W=1.25E-06 $X=7945 $Y=15880 $D=1
M285 10 47 VDD VDD P12LL L=6E-08 W=1E-06 $X=8235 $Y=1195 $D=1
M286 50 45 VDD VDD P12LL L=6E-08 W=1E-06 $X=8235 $Y=3025 $D=1
M287 48 49 VDD VDD P12LL L=6E-08 W=4E-07 $X=8235 $Y=9125 $D=1
M288 FCKX[5] 49 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=8235 $Y=12320 $D=1
M289 FCKX[5] 48 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=8235 $Y=15880 $D=1
M290 49 48 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=8325 $Y=8285 $D=1
M291 49 CLK 50 VDD P12LL L=6E-08 W=5E-07 $X=8395 $Y=7170 $D=1
M292 VDD 47 10 VDD P12LL L=6E-08 W=1E-06 $X=8525 $Y=1195 $D=1
M293 VDD 53 50 VDD P12LL L=6E-08 W=1E-06 $X=8525 $Y=3025 $D=1
M294 VDD 49 48 VDD P12LL L=6E-08 W=4E-07 $X=8525 $Y=9125 $D=1
M295 WLCKX 49 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=8525 $Y=12320 $D=1
M296 VDD 48 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=8525 $Y=15880 $D=1
M297 50 CLK 49 VDD P12LL L=6E-08 W=5E-07 $X=8675 $Y=7170 $D=1
M298 53 10 VDD VDD P12LL L=6E-08 W=1E-06 $X=8815 $Y=1195 $D=1
M299 50 5 VDD VDD P12LL L=6E-08 W=1E-06 $X=8815 $Y=3025 $D=1
M300 48 49 VDD VDD P12LL L=6E-08 W=4E-07 $X=8815 $Y=9125 $D=1
M301 FCKX[5] 49 WLCKX VDD P12LL L=6E-08 W=1.25E-06 $X=8815 $Y=12320 $D=1
M302 FCKX[5] 48 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=8815 $Y=15880 $D=1
M303 49 CLK 50 VDD P12LL L=6E-08 W=5E-07 $X=8945 $Y=7170 $D=1
M304 VDD 10 53 VDD P12LL L=6E-08 W=1E-06 $X=9105 $Y=1195 $D=1
M305 VDD 49 48 VDD P12LL L=6E-08 W=4E-07 $X=9105 $Y=9125 $D=1
M306 WLCKX 49 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=9105 $Y=12320 $D=1
M307 VDD 48 FCKX[5] VDD P12LL L=6E-08 W=1.25E-06 $X=9105 $Y=15880 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLSTRAP_B                                                            *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBLSTRAP_B VDD VSS BL BLX
*.NOPIN VSS
*.PININFO BL:B BLX:B 
MTA1 BLX VSS NET7 VSS RFNPGBHVT W=0.12U L=0.09U M=1
MTA0 BL VSS NET4 VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTD1 NET11 VSS VSS VSS RFNPDHVT W=0.46U L=0.07U M=1
MTL1 VDD VSS NET12 VDD RFPLHVT W=0.095U L=0.07U M=1
.ENDS qspi_data_info_32_memBLSTRAP_B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL                                                          *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL VDD VSS BA BB BXA BXB WLA
*.NOPIN VSS
*.PININFO BA:B BB:B BXA:B BXB:B WLA:I 
MTD0 VSS BCN BC VSS RFNPDHVT W=0.46U L=0.07U M=1
MN2 BXB VSS BCN VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTA1 BXA WLA BCN VSS RFNPGBHVT W=0.12U L=0.09U M=1
MN1 BC VSS BB VSS RFNPGBHVT W=0.12U L=0.09U M=1
MTA0 BC WLA BA VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTD1 BCN BC VSS VSS RFNPDHVT W=0.46U L=0.07U M=1
MTL1 VDD BC BCN VDD RFPLHVT W=0.095U L=0.07U M=1
MTL0 BC BCN VDD VDD RFPLHVT W=0.095U L=0.07U M=1
.ENDS qspi_data_info_32_memTP_EDGECELL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL8A                                                        *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL8A VDD VSS BA0 BA7 BXA0 BXA7 WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BA0:B BA7:B BXA0:B BXA7:B WLA[7]:I WLA[6]:I WLA[5]:I WLA[4]:I
*.PININFO WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS NET0105 NET19 NET20 NET050 WLA[4] qspi_data_info_32_memTP_EDGECELL
XI6 VDD VSS NET095 NET19 NET076 NET050 WLA[5] qspi_data_info_32_memTP_EDGECELL
XI5 VDD VSS BA7 NET036 BXA7 NET040 WLA[7] qspi_data_info_32_memTP_EDGECELL
XI4 VDD VSS NET095 NET036 NET076 NET040 WLA[6] qspi_data_info_32_memTP_EDGECELL
XI3 VDD VSS NET0115 NET056 NET24 NET055 WLA[2] qspi_data_info_32_memTP_EDGECELL
XI2 VDD VSS NET0105 NET056 NET20 NET055 WLA[3] qspi_data_info_32_memTP_EDGECELL
XI1 VDD VSS NET0115 NET091 NET24 NET030 WLA[1] qspi_data_info_32_memTP_EDGECELL
XI0 VDD VSS BA0 NET091 BXA0 NET030 WLA[0] qspi_data_info_32_memTP_EDGECELL
.ENDS qspi_data_info_32_memTP_EDGECELL8A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL34B                                                       *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL34B VDD VSS RWL[0] RWL[1] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO RWL[0]:I RWL[1]:I WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I
*.PININFO WLA[26]:I WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I
*.PININFO WLA[19]:I WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I
*.PININFO WLA[12]:I WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I
*.PININFO WLA[5]:I WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI4 VDD VSS NET33 NET32 qspi_data_info_32_memBLSTRAP_B
XI5 VDD VSS NET035 NET034 qspi_data_info_32_memBLSTRAP_B
XI6 VDD VSS NET028 NET057 NET027 NET056 RWL[1] qspi_data_info_32_memTP_EDGECELL
XI7 VDD VSS NET035 NET057 NET034 NET056 RWL[0] qspi_data_info_32_memTP_EDGECELL
XI2 VDD VSS NET028 NET14 NET027 NET13 WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1]
+WLA[0] qspi_data_info_32_memTP_EDGECELL8A
XI3 VDD VSS NET043 NET14 NET042 NET13 WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] qspi_data_info_32_memTP_EDGECELL8A
XI1 VDD VSS NET043 NET28 NET042 NET27 WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] qspi_data_info_32_memTP_EDGECELL8A
XI0 VDD VSS NET33 NET28 NET32 NET27 WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] qspi_data_info_32_memTP_EDGECELL8A
.ENDS qspi_data_info_32_memTP_EDGECELL34B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLSTRAP_A                                                            *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBLSTRAP_A VDD VSS BL BLX
*.NOPIN VSS
*.PININFO BL:B BLX:B 
MTA1 BLX VSS NET7 VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTA0 BL VSS NET4 VSS RFNPGBHVT W=0.12U L=0.09U M=1
MTD1 NET11 VSS VSS VSS RFNPDHVT W=0.46U L=0.07U M=1
MTL1 VDD VSS NET12 VDD RFPLHVT W=0.095U L=0.07U M=1
.ENDS qspi_data_info_32_memBLSTRAP_A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL8B                                                        *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL8B VDD VSS BB0 BB7 BXB0 BXB7 WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BB0:B BB7:B BXB0:B BXB7:B WLA[7]:I WLA[6]:I WLA[5]:I WLA[4]:I
*.PININFO WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS NET095 NET19 NET20 NET050 WLA[4] qspi_data_info_32_memTP_EDGECELL
XI6 VDD VSS NET095 NET057 NET20 NET034 WLA[5] qspi_data_info_32_memTP_EDGECELL
XI5 VDD VSS NET054 BB7 NET053 BXB7 WLA[7] qspi_data_info_32_memTP_EDGECELL
XI4 VDD VSS NET054 NET057 NET053 NET034 WLA[6] qspi_data_info_32_memTP_EDGECELL
XI3 VDD VSS NET0115 NET091 NET24 NET055 WLA[2] qspi_data_info_32_memTP_EDGECELL
XI2 VDD VSS NET0115 NET19 NET24 NET050 WLA[3] qspi_data_info_32_memTP_EDGECELL
XI1 VDD VSS NET074 NET091 NET073 NET055 WLA[1] qspi_data_info_32_memTP_EDGECELL
XI0 VDD VSS NET074 BB0 NET073 BXB0 WLA[0] qspi_data_info_32_memTP_EDGECELL
.ENDS qspi_data_info_32_memTP_EDGECELL8B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL32A                                                       *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL32A VDD VSS WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25]
+WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I WLA[26]:I WLA[25]:I
*.PININFO WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I WLA[19]:I WLA[18]:I
*.PININFO WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I WLA[12]:I WLA[11]:I
*.PININFO WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I WLA[5]:I WLA[4]:I
*.PININFO WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI4 VDD VSS NET57 NET56 qspi_data_info_32_memBLSTRAP_A
XI5 VDD VSS NET62 NET045 qspi_data_info_32_memBLSTRAP_A
XI2 VDD VSS NET62 NET42 NET045 NET61 WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] qspi_data_info_32_memTP_EDGECELL8B
XI3 VDD VSS NET47 NET42 NET51 NET61 WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] qspi_data_info_32_memTP_EDGECELL8B
XI1 VDD VSS NET47 NET034 NET51 NET033 WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] qspi_data_info_32_memTP_EDGECELL8B
XI0 VDD VSS NET57 NET034 NET56 NET033 WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1]
+WLA[0] qspi_data_info_32_memTP_EDGECELL8B
.ENDS qspi_data_info_32_memTP_EDGECELL32A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_EDGECELL64AB                                                     *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_EDGECELL64AB VDD VSS RWL[0] RWL[1] WLA[63] WLA[62] 
+WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] 
+WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] 
+WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] 
+WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] 
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] 
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] 
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
XI3 VDD VSS RWL[0] RWL[1] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25]
+WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16]
+WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6]
+WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] qspi_data_info_32_memTP_EDGECELL34B
XI8_2 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] 
+WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] 
+WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] 
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] 
+qspi_data_info_32_memTP_EDGECELL32A
.ENDS qspi_data_info_32_memTP_EDGECELL64AB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL                                                              *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL VDD VSS BA BB BXA BXB WLA WLB
*.NOPIN VSS
*.PININFO BA:B BB:B BXA:B BXB:B WLA:I WLB:I 
MTD0 VSS BCN BC VSS RFNPDHVT W=0.46U L=0.07U M=1
MN2 BXB WLB BCN VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTA1 BXA WLA BCN VSS RFNPGBHVT W=0.12U L=0.09U M=1
MN1 BC WLB BB VSS RFNPGBHVT W=0.12U L=0.09U M=1
MTA0 BC WLA BA VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTD1 BCN BC VSS VSS RFNPDHVT W=0.46U L=0.07U M=1
MTL1 VDD BC BCN VDD RFPLHVT W=0.095U L=0.07U M=1
MTL0 BC BCN VDD VDD RFPLHVT W=0.095U L=0.07U M=1
.ENDS qspi_data_info_32_memBITCELL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL2X2                                                           *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL2X2 VDD VSS BA[1] BA[0] BB[1] BB[0] BXA[1] BXA[0] BXB[1] BXB[0] WLA[0]
+WLA[1] WLB[0] WLB[1]
*.NOPIN VSS
*.PININFO BA[1]:B BA[0]:B BB[1]:B BB[0]:B BXA[1]:B BXA[0]:B BXB[1]:B BXB[0]:B
*.PININFO WLA[0]:I WLA[1]:I WLB[0]:I WLB[1]:I 
XI3 VDD VSS BA[1] BB[1] BXA[1] BXB[1] WLA[1] WLB[1] qspi_data_info_32_memBITCELL
XI2 VDD VSS BA[1] BB[1] BXA[1] BXB[1] WLA[0] WLB[0] qspi_data_info_32_memBITCELL
XI1 VDD VSS BA[0] BB[0] BXA[0] BXB[0] WLA[1] WLB[1] qspi_data_info_32_memBITCELL
XI0 VDD VSS BA[0] BB[0] BXA[0] BXB[0] WLA[0] WLB[0] qspi_data_info_32_memBITCELL
.ENDS qspi_data_info_32_memBITCELL2X2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL32X1A                                                         *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL32X1A VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25]
+WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI3_1 VDD VSS BLB[1] BLXB[1] qspi_data_info_32_memBLSTRAP_A
XI3_0 VDD VSS BLB[0] BLXB[0] qspi_data_info_32_memBLSTRAP_A
XI1_1 VDD VSS BLB[1] BLXB[1] qspi_data_info_32_memBLSTRAP_A
XI1_0 VDD VSS BLB[0] BLXB[0] qspi_data_info_32_memBLSTRAP_A
XI0_15 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[31] WLA[30] WLB[31] WLB[30] qspi_data_info_32_memBITCELLB2X1
XI0_14 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[29] WLA[28] WLB[29] WLB[28] qspi_data_info_32_memBITCELLB2X1
XI0_13 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[27] WLA[26] WLB[27] WLB[26] qspi_data_info_32_memBITCELLB2X1
XI0_12 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[25] WLA[24] WLB[25] WLB[24] qspi_data_info_32_memBITCELLB2X1
XI0_11 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[23] WLA[22] WLB[23] WLB[22] qspi_data_info_32_memBITCELLB2X1
XI0_10 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[21] WLA[20] WLB[21] WLB[20] qspi_data_info_32_memBITCELLB2X1
XI0_9 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[19] WLA[18] WLB[19] WLB[18] qspi_data_info_32_memBITCELLB2X1
XI0_8 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[17] WLA[16] WLB[17] WLB[16] qspi_data_info_32_memBITCELLB2X1
XI0_7 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[15] WLA[14] WLB[15] WLB[14] qspi_data_info_32_memBITCELLB2X1
XI0_6 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[13] WLA[12] WLB[13] WLB[12] qspi_data_info_32_memBITCELLB2X1
XI0_5 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[11] WLA[10] WLB[11] WLB[10] qspi_data_info_32_memBITCELLB2X1
XI0_4 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[9] WLA[8] WLB[9] WLB[8] qspi_data_info_32_memBITCELLB2X1
XI0_3 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[7] WLA[6] WLB[7] WLB[6] qspi_data_info_32_memBITCELLB2X1
XI0_2 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[5] WLA[4] WLB[5] WLB[4] qspi_data_info_32_memBITCELLB2X1
XI0_1 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[3] WLA[2] WLB[3] WLB[2] qspi_data_info_32_memBITCELLB2X1
XI0_0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[1] WLA[0] WLB[1] WLB[0] qspi_data_info_32_memBITCELLB2X1
.ENDS qspi_data_info_32_memBITCELL32X1A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL2X1_RD                                                        *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL2X1_RD VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[0] WLA[1] WLB[0] WLB[1]
XI0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] WLA[0] WLA[1]
+WLB[0] WLB[1] qspi_data_info_32_memBITCELL2X2
.ENDS qspi_data_info_32_memBITCELL2X1_RD


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL34X1B                                                         *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL34X1B VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[31] WLB[30] WLB[29]
+WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11]
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI3_1 VDD VSS BLA[1] BLXA[1] qspi_data_info_32_memBLSTRAP_B
XI3_0 VDD VSS BLA[0] BLXA[0] qspi_data_info_32_memBLSTRAP_B
XI1_1 VDD VSS BLA[1] BLXA[1] qspi_data_info_32_memBLSTRAP_B
XI1_0 VDD VSS BLA[0] BLXA[0] qspi_data_info_32_memBLSTRAP_B
XI4 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1] qspi_data_info_32_memBITCELL2X1_RD
XI0_15 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[31] WLA[30] WLB[31] WLB[30] qspi_data_info_32_memBITCELLB2X1
XI0_14 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[29] WLA[28] WLB[29] WLB[28] qspi_data_info_32_memBITCELLB2X1
XI0_13 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[27] WLA[26] WLB[27] WLB[26] qspi_data_info_32_memBITCELLB2X1
XI0_12 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[25] WLA[24] WLB[25] WLB[24] qspi_data_info_32_memBITCELLB2X1
XI0_11 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[23] WLA[22] WLB[23] WLB[22] qspi_data_info_32_memBITCELLB2X1
XI0_10 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[21] WLA[20] WLB[21] WLB[20] qspi_data_info_32_memBITCELLB2X1
XI0_9 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[19] WLA[18] WLB[19] WLB[18] qspi_data_info_32_memBITCELLB2X1
XI0_8 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[17] WLA[16] WLB[17] WLB[16] qspi_data_info_32_memBITCELLB2X1
XI0_7 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[15] WLA[14] WLB[15] WLB[14] qspi_data_info_32_memBITCELLB2X1
XI0_6 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[13] WLA[12] WLB[13] WLB[12] qspi_data_info_32_memBITCELLB2X1
XI0_5 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[11] WLA[10] WLB[11] WLB[10] qspi_data_info_32_memBITCELLB2X1
XI0_4 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[9] WLA[8] WLB[9] WLB[8] qspi_data_info_32_memBITCELLB2X1
XI0_3 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[7] WLA[6] WLB[7] WLB[6] qspi_data_info_32_memBITCELLB2X1
XI0_2 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[5] WLA[4] WLB[5] WLB[4] qspi_data_info_32_memBITCELLB2X1
XI0_1 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[3] WLA[2] WLB[3] WLB[2] qspi_data_info_32_memBITCELLB2X1
XI0_0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[1] WLA[0] WLB[1] WLB[0] qspi_data_info_32_memBITCELLB2X1
.ENDS qspi_data_info_32_memBITCELL34X1B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELL32X1B                                                         *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELL32X1B VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22]
+WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13]
+WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25]
+WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16]
+WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] WLB[6]
+WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
XI3_1 VDD VSS BLA[1] BLXA[1] qspi_data_info_32_memBLSTRAP_B
XI3_0 VDD VSS BLA[0] BLXA[0] qspi_data_info_32_memBLSTRAP_B
XI1_1 VDD VSS BLA[1] BLXA[1] qspi_data_info_32_memBLSTRAP_B
XI1_0 VDD VSS BLA[0] BLXA[0] qspi_data_info_32_memBLSTRAP_B
XI0_15 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[31] WLA[30] WLB[31] WLB[30] qspi_data_info_32_memBITCELLB2X1
XI0_14 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[29] WLA[28] WLB[29] WLB[28] qspi_data_info_32_memBITCELLB2X1
XI0_13 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[27] WLA[26] WLB[27] WLB[26] qspi_data_info_32_memBITCELLB2X1
XI0_12 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[25] WLA[24] WLB[25] WLB[24] qspi_data_info_32_memBITCELLB2X1
XI0_11 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[23] WLA[22] WLB[23] WLB[22] qspi_data_info_32_memBITCELLB2X1
XI0_10 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[21] WLA[20] WLB[21] WLB[20] qspi_data_info_32_memBITCELLB2X1
XI0_9 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[19] WLA[18] WLB[19] WLB[18] qspi_data_info_32_memBITCELLB2X1
XI0_8 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[17] WLA[16] WLB[17] WLB[16] qspi_data_info_32_memBITCELLB2X1
XI0_7 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[15] WLA[14] WLB[15] WLB[14] qspi_data_info_32_memBITCELLB2X1
XI0_6 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[13] WLA[12] WLB[13] WLB[12] qspi_data_info_32_memBITCELLB2X1
XI0_5 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[11] WLA[10] WLB[11] WLB[10] qspi_data_info_32_memBITCELLB2X1
XI0_4 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[9] WLA[8] WLB[9] WLB[8] qspi_data_info_32_memBITCELLB2X1
XI0_3 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[7] WLA[6] WLB[7] WLB[6] qspi_data_info_32_memBITCELLB2X1
XI0_2 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[5] WLA[4] WLB[5] WLB[4] qspi_data_info_32_memBITCELLB2X1
XI0_1 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[3] WLA[2] WLB[3] WLB[2] qspi_data_info_32_memBITCELLB2X1
XI0_0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[1] WLA[0] WLB[1] WLB[0] qspi_data_info_32_memBITCELLB2X1
.ENDS qspi_data_info_32_memBITCELL32X1B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: ARRAY64X1                                                           *
*******************************************************************************
.SUBCKT qspi_data_info_32_memARRAY64X1 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] 
+WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] 
+WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] 
+WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] 
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] 
+WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] 
+WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8] WLB[7] 
+WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
XI4 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24]
+WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15]
+WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5]
+WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27]
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18]
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] WLB[8]
+WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] qspi_data_info_32_memBITCELL34X1B
XI5_1 VDD VSS BLXA[1] BLXA[0] BLXB[1] BLXB[0] BLA[1] BLA[0] BLB[1] BLB[0]
+WLA[63] WLA[62] WLA[61] WLA[60] WLA[59] 
+WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] 
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] 
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] 
+WLB[63] WLB[62] WLB[61] WLB[60] WLB[59] 
+WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50] 
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] 
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] 
+qspi_data_info_32_memBITCELL32X1A
.ENDS qspi_data_info_32_memARRAY64X1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YMX1R                                                              *
*******************************************************************************
.SUBCKT qspi_data_info_32_memYMX1R VDD VSS DB[1] DB[0] DBX[1] DBX[0] DOUT[1] DOUT[0] CK1 CK4

M0 34 14 VSS VSS N12LL L=6E-08 W=1E-06 $X=485 $Y=12550 $D=0
M1 27 11 34 VSS N12LL L=6E-08 W=1E-06 $X=485 $Y=12790 $D=0
M2 8 13 27 VSS N12LL L=1.2E-07 W=1E-06 $X=490 $Y=13280 $D=0
M3 VSS 23 10 VSS N12LL L=6E-08 W=5E-07 $X=515 $Y=6185 $D=0
M4 VSS CK1 22 VSS N12LL L=6E-08 W=4E-07 $X=530 $Y=4905 $D=0
M5 35 8 24 VSS N12LL L=6E-08 W=1E-06 $X=705 $Y=10995 $D=0
M6 36 CK1 VSS VSS N12LL L=6E-08 W=4E-07 $X=805 $Y=6285 $D=0
M7 11 22 VSS VSS N12LL L=6E-08 W=4E-07 $X=810 $Y=4905 $D=0
M8 27 13 8 VSS N12LL L=1.2E-07 W=1E-06 $X=880 $Y=13280 $D=0
M9 VSS 26 35 VSS N12LL L=6E-08 W=1E-06 $X=960 $Y=10995 $D=0
M10 23 CK4 36 VSS N12LL L=6E-08 W=4E-07 $X=1035 $Y=6285 $D=0
M11 37 24 VSS VSS N12LL L=6E-08 W=1E-06 $X=1250 $Y=10995 $D=0
M12 13 8 27 VSS N12LL L=1.2E-07 W=1E-06 $X=1270 $Y=13280 $D=0
M13 26 13 37 VSS N12LL L=6E-08 W=1E-06 $X=1505 $Y=10995 $D=0
M14 VSS CK4 25 VSS N12LL L=6E-08 W=4E-07 $X=1555 $Y=4910 $D=0
M15 27 8 13 VSS N12LL L=1.2E-07 W=1E-06 $X=1660 $Y=13280 $D=0
M16 DOUT[0] 24 VSS VSS N12LL L=6E-08 W=7E-07 $X=1805 $Y=5995 $D=0
M17 14 25 VSS VSS N12LL L=6E-08 W=4E-07 $X=1825 $Y=4910 $D=0
M18 VSS 25 14 VSS N12LL L=6E-08 W=4E-07 $X=2095 $Y=4910 $D=0
M19 VSS 24 DOUT[0] VSS N12LL L=6E-08 W=7E-07 $X=2095 $Y=5995 $D=0
M20 16 28 VSS VSS N12LL L=6E-08 W=4E-07 $X=2385 $Y=4910 $D=0
M21 DOUT[1] 31 VSS VSS N12LL L=6E-08 W=7E-07 $X=2385 $Y=5995 $D=0
M22 VSS 28 16 VSS N12LL L=6E-08 W=4E-07 $X=2655 $Y=4910 $D=0
M23 VSS 31 DOUT[1] VSS N12LL L=6E-08 W=7E-07 $X=2675 $Y=5995 $D=0
M24 15 19 33 VSS N12LL L=1.2E-07 W=1E-06 $X=2760 $Y=13280 $D=0
M25 28 CK4 VSS VSS N12LL L=6E-08 W=4E-07 $X=2925 $Y=4910 $D=0
M26 38 15 29 VSS N12LL L=6E-08 W=1E-06 $X=2975 $Y=10995 $D=0
M27 39 16 VSS VSS N12LL L=6E-08 W=1E-06 $X=3055 $Y=12550 $D=0
M28 33 17 39 VSS N12LL L=6E-08 W=1E-06 $X=3055 $Y=12790 $D=0
M29 33 19 15 VSS N12LL L=1.2E-07 W=1E-06 $X=3150 $Y=13280 $D=0
M30 VSS 31 38 VSS N12LL L=6E-08 W=1E-06 $X=3230 $Y=10995 $D=0
M31 40 CK4 30 VSS N12LL L=6E-08 W=4E-07 $X=3445 $Y=6285 $D=0
M32 41 29 VSS VSS N12LL L=6E-08 W=1E-06 $X=3520 $Y=10995 $D=0
M33 19 15 33 VSS N12LL L=1.2E-07 W=1E-06 $X=3540 $Y=13280 $D=0
M34 VSS 32 17 VSS N12LL L=6E-08 W=4E-07 $X=3670 $Y=4905 $D=0
M35 VSS CK1 40 VSS N12LL L=6E-08 W=4E-07 $X=3675 $Y=6285 $D=0
M36 31 19 41 VSS N12LL L=6E-08 W=1E-06 $X=3775 $Y=10995 $D=0
M37 33 15 19 VSS N12LL L=1.2E-07 W=1E-06 $X=3930 $Y=13280 $D=0
M38 32 CK1 VSS VSS N12LL L=6E-08 W=4E-07 $X=3950 $Y=4905 $D=0
M39 20 30 VSS VSS N12LL L=6E-08 W=5E-07 $X=3965 $Y=6185 $D=0
M40 8 13 VDD VDD P12LL L=1.2E-07 W=4E-07 $X=490 $Y=15180 $D=1
M41 DB[0] 10 8 VDD P12LL L=6E-08 W=5E-07 $X=500 $Y=16365 $D=1
M42 VDD 23 10 VDD P12LL L=6E-08 W=1E-06 $X=515 $Y=7495 $D=1
M43 VDD CK1 22 VDD P12LL L=6E-08 W=4E-07 $X=530 $Y=3615 $D=1
M44 24 8 VDD VDD P12LL L=6E-08 W=1E-06 $X=670 $Y=9170 $D=1
M45 8 10 DB[0] VDD P12LL L=6E-08 W=5E-07 $X=790 $Y=16365 $D=1
M46 23 CK1 VDD VDD P12LL L=6E-08 W=4E-07 $X=805 $Y=7495 $D=1
M47 11 22 VDD VDD P12LL L=6E-08 W=4E-07 $X=810 $Y=3615 $D=1
M48 DB[0] 14 VDD VDD P12LL L=6E-08 W=1E-06 $X=815 $Y=17430 $D=1
M49 VDD 13 8 VDD P12LL L=1.2E-07 W=4E-07 $X=880 $Y=15180 $D=1
M50 VDD 26 24 VDD P12LL L=6E-08 W=1E-06 $X=960 $Y=9170 $D=1
M51 VDD CK4 23 VDD P12LL L=6E-08 W=4E-07 $X=1095 $Y=7495 $D=1
M52 DBX[0] 14 DB[0] VDD P12LL L=6E-08 W=1E-06 $X=1105 $Y=17430 $D=1
M53 26 24 VDD VDD P12LL L=6E-08 W=1E-06 $X=1250 $Y=9170 $D=1
M54 13 8 VDD VDD P12LL L=1.2E-07 W=4E-07 $X=1270 $Y=15180 $D=1
M55 VDD 14 DBX[0] VDD P12LL L=6E-08 W=1E-06 $X=1395 $Y=17430 $D=1
M56 DBX[0] 10 13 VDD P12LL L=6E-08 W=5E-07 $X=1420 $Y=16365 $D=1
M57 VDD 13 26 VDD P12LL L=6E-08 W=1E-06 $X=1540 $Y=9170 $D=1
M58 VDD CK4 25 VDD P12LL L=6E-08 W=8E-07 $X=1555 $Y=3285 $D=1
M59 VDD 8 13 VDD P12LL L=1.2E-07 W=4E-07 $X=1660 $Y=15180 $D=1
M60 13 10 DBX[0] VDD P12LL L=6E-08 W=5E-07 $X=1710 $Y=16365 $D=1
M61 DOUT[0] 24 VDD VDD P12LL L=6E-08 W=1.2E-06 $X=1805 $Y=7495 $D=1
M62 14 25 VDD VDD P12LL L=6E-08 W=8E-07 $X=1825 $Y=3285 $D=1
M63 VDD 25 14 VDD P12LL L=6E-08 W=8E-07 $X=2095 $Y=3285 $D=1
M64 VDD 24 DOUT[0] VDD P12LL L=6E-08 W=1.2E-06 $X=2095 $Y=7495 $D=1
M65 16 28 VDD VDD P12LL L=6E-08 W=8E-07 $X=2385 $Y=3285 $D=1
M66 DOUT[1] 31 VDD VDD P12LL L=6E-08 W=1.2E-06 $X=2385 $Y=7495 $D=1
M67 VDD 28 16 VDD P12LL L=6E-08 W=8E-07 $X=2655 $Y=3285 $D=1
M68 VDD 31 DOUT[1] VDD P12LL L=6E-08 W=1.2E-06 $X=2675 $Y=7495 $D=1
M69 15 19 VDD VDD P12LL L=1.2E-07 W=4E-07 $X=2760 $Y=15180 $D=1
M70 DBX[1] 20 15 VDD P12LL L=6E-08 W=5E-07 $X=2770 $Y=16365 $D=1
M71 28 CK4 VDD VDD P12LL L=6E-08 W=8E-07 $X=2925 $Y=3285 $D=1
M72 29 15 VDD VDD P12LL L=6E-08 W=1E-06 $X=2940 $Y=9170 $D=1
M73 15 20 DBX[1] VDD P12LL L=6E-08 W=5E-07 $X=3060 $Y=16365 $D=1
M74 DBX[1] 16 VDD VDD P12LL L=6E-08 W=1E-06 $X=3085 $Y=17430 $D=1
M75 VDD 19 15 VDD P12LL L=1.2E-07 W=4E-07 $X=3150 $Y=15180 $D=1
M76 VDD 31 29 VDD P12LL L=6E-08 W=1E-06 $X=3230 $Y=9170 $D=1
M77 DB[1] 16 DBX[1] VDD P12LL L=6E-08 W=1E-06 $X=3375 $Y=17430 $D=1
M78 30 CK4 VDD VDD P12LL L=6E-08 W=4E-07 $X=3385 $Y=7495 $D=1
M79 31 29 VDD VDD P12LL L=6E-08 W=1E-06 $X=3520 $Y=9170 $D=1
M80 19 15 VDD VDD P12LL L=1.2E-07 W=4E-07 $X=3540 $Y=15180 $D=1
M81 VDD 16 DB[1] VDD P12LL L=6E-08 W=1E-06 $X=3665 $Y=17430 $D=1
M82 VDD 32 17 VDD P12LL L=6E-08 W=4E-07 $X=3670 $Y=3615 $D=1
M83 VDD CK1 30 VDD P12LL L=6E-08 W=4E-07 $X=3675 $Y=7495 $D=1
M84 DB[1] 20 19 VDD P12LL L=6E-08 W=5E-07 $X=3690 $Y=16365 $D=1
M85 VDD 19 31 VDD P12LL L=6E-08 W=1E-06 $X=3810 $Y=9170 $D=1
M86 VDD 15 19 VDD P12LL L=1.2E-07 W=4E-07 $X=3930 $Y=15180 $D=1
M87 32 CK1 VDD VDD P12LL L=6E-08 W=4E-07 $X=3950 $Y=3615 $D=1
M88 20 30 VDD VDD P12LL L=6E-08 W=1E-06 $X=3965 $Y=7495 $D=1
M89 19 20 DB[1] VDD P12LL L=6E-08 W=5E-07 $X=3980 $Y=16365 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YMX1W                                                              *
*******************************************************************************
.SUBCKT qspi_data_info_32_memYMX1W VDD VSS BLW[1] BLW[0] BLXW[1] BLXW[0] BWEN[1] BWEN[0] CTRCLKW CTRCLKWX
+DATA[1] DATA[0] INTCLKX

M0 45 VDD VSS VSS N12LL L=4E-07 W=4E-07 $X=145 $Y=5385 $D=0
M1 44 9 VSS VSS N12LL L=6E-08 W=1.2E-07 $X=170 $Y=12935 $D=0
M2 47 VDD VSS VSS N12LL L=4E-07 W=4E-07 $X=375 $Y=1050 $D=0
M3 32 CTRCLKW 44 VSS N12LL L=6E-08 W=1.2E-07 $X=450 $Y=12935 $D=0
M4 BLXW[0] 9 37 VSS N12LL L=6E-08 W=1E-06 $X=560 $Y=17935 $D=0
M5 9 32 VSS VSS N12LL L=6E-08 W=1E-06 $X=575 $Y=14270 $D=0
M6 46 13 10 VSS N12LL L=6E-08 W=1.2E-06 $X=680 $Y=7070 $D=0
M7 33 12 45 VSS N12LL L=3E-07 W=4E-07 $X=745 $Y=5385 $D=0
M8 10 CTRCLKWX 32 VSS N12LL L=6E-08 W=1.2E-06 $X=790 $Y=12465 $D=0
M9 37 9 BLXW[0] VSS N12LL L=6E-08 W=1E-06 $X=830 $Y=17935 $D=0
M10 VSS 32 9 VSS N12LL L=6E-08 W=1E-06 $X=865 $Y=14270 $D=0
M11 VSS 33 46 VSS N12LL L=6E-08 W=1.2E-06 $X=960 $Y=7070 $D=0
M12 17 DATA[0] 47 VSS N12LL L=3E-07 W=4E-07 $X=975 $Y=1050 $D=0
M13 VSS 36 37 VSS N12LL L=6E-08 W=1E-06 $X=1100 $Y=17935 $D=0
M14 18 35 VSS VSS N12LL L=6E-08 W=1E-06 $X=1155 $Y=14270 $D=0
M15 48 33 VSS VSS N12LL L=6E-08 W=1.2E-06 $X=1250 $Y=7070 $D=0
M16 37 36 VSS VSS N12LL L=6E-08 W=1E-06 $X=1370 $Y=17935 $D=0
M17 35 CTRCLKWX 15 VSS N12LL L=6E-08 W=1.2E-06 $X=1420 $Y=12465 $D=0
M18 VSS 35 18 VSS N12LL L=6E-08 W=1E-06 $X=1445 $Y=14270 $D=0
M19 VSS 34 12 VSS N12LL L=6E-08 W=6E-07 $X=1480 $Y=5975 $D=0
M20 15 17 48 VSS N12LL L=6E-08 W=1.2E-06 $X=1530 $Y=7070 $D=0
M21 BLW[0] 18 37 VSS N12LL L=6E-08 W=1E-06 $X=1640 $Y=17935 $D=0
M22 13 17 VSS VSS N12LL L=6E-08 W=4E-07 $X=1760 $Y=5975 $D=0
M23 49 CTRCLKW 35 VSS N12LL L=6E-08 W=1.2E-07 $X=1760 $Y=12935 $D=0
M24 VSS VSS DATA[0] VSS N12LL L=6E-08 W=2E-07 $X=1865 $Y=1065 $D=0
M25 37 18 BLW[0] VSS N12LL L=6E-08 W=1E-06 $X=1910 $Y=17935 $D=0
M26 VSS 18 49 VSS N12LL L=6E-08 W=1.2E-07 $X=2040 $Y=12935 $D=0
M27 VSS INTCLKX 36 VSS N12LL L=6E-08 W=6E-07 $X=2095 $Y=14565 $D=0
M28 38 INTCLKX VSS VSS N12LL L=6E-08 W=6E-07 $X=2385 $Y=14565 $D=0
M29 50 22 VSS VSS N12LL L=6E-08 W=1.2E-07 $X=2440 $Y=12935 $D=0
M30 BLW[1] 22 43 VSS N12LL L=6E-08 W=1E-06 $X=2570 $Y=17935 $D=0
M31 DATA[1] VSS VSS VSS N12LL L=6E-08 W=2E-07 $X=2615 $Y=1065 $D=0
M32 VSS 20 29 VSS N12LL L=6E-08 W=4E-07 $X=2720 $Y=5975 $D=0
M33 39 CTRCLKW 50 VSS N12LL L=6E-08 W=1.2E-07 $X=2720 $Y=12935 $D=0
M34 43 22 BLW[1] VSS N12LL L=6E-08 W=1E-06 $X=2840 $Y=17935 $D=0
M35 51 20 24 VSS N12LL L=6E-08 W=1.2E-06 $X=2950 $Y=7070 $D=0
M36 26 40 VSS VSS N12LL L=6E-08 W=6E-07 $X=3000 $Y=5975 $D=0
M37 22 39 VSS VSS N12LL L=6E-08 W=1E-06 $X=3035 $Y=14270 $D=0
M38 24 CTRCLKWX 39 VSS N12LL L=6E-08 W=1.2E-06 $X=3060 $Y=12465 $D=0
M39 VSS 38 43 VSS N12LL L=6E-08 W=1E-06 $X=3110 $Y=17935 $D=0
M40 VSS 41 51 VSS N12LL L=6E-08 W=1.2E-06 $X=3230 $Y=7070 $D=0
M41 52 DATA[1] 20 VSS N12LL L=3E-07 W=4E-07 $X=3265 $Y=1050 $D=0
M42 VSS 39 22 VSS N12LL L=6E-08 W=1E-06 $X=3325 $Y=14270 $D=0
M43 43 38 VSS VSS N12LL L=6E-08 W=1E-06 $X=3380 $Y=17935 $D=0
M44 54 26 41 VSS N12LL L=3E-07 W=4E-07 $X=3495 $Y=5385 $D=0
M45 53 41 VSS VSS N12LL L=6E-08 W=1.2E-06 $X=3520 $Y=7070 $D=0
M46 31 42 VSS VSS N12LL L=6E-08 W=1E-06 $X=3615 $Y=14270 $D=0
M47 BLXW[1] 31 43 VSS N12LL L=6E-08 W=1E-06 $X=3650 $Y=17935 $D=0
M48 42 CTRCLKWX 27 VSS N12LL L=6E-08 W=1.2E-06 $X=3690 $Y=12465 $D=0
M49 VSS VDD 52 VSS N12LL L=4E-07 W=4E-07 $X=3765 $Y=1050 $D=0
M50 27 29 53 VSS N12LL L=6E-08 W=1.2E-06 $X=3800 $Y=7070 $D=0
M51 VSS 42 31 VSS N12LL L=6E-08 W=1E-06 $X=3905 $Y=14270 $D=0
M52 43 31 BLXW[1] VSS N12LL L=6E-08 W=1E-06 $X=3920 $Y=17935 $D=0
M53 VSS VDD 54 VSS N12LL L=4E-07 W=4E-07 $X=3995 $Y=5385 $D=0
M54 55 CTRCLKW 42 VSS N12LL L=6E-08 W=1.2E-07 $X=4030 $Y=12935 $D=0
M55 VSS 31 55 VSS N12LL L=6E-08 W=1.2E-07 $X=4310 $Y=12935 $D=0
M56 57 VSS VDD VDD P12LL L=2E-07 W=4E-07 $X=140 $Y=4300 $D=1
M57 56 9 VDD VDD P12LL L=6E-08 W=1.2E-07 $X=170 $Y=11815 $D=1
M58 32 CTRCLKWX 56 VDD P12LL L=6E-08 W=1.2E-07 $X=450 $Y=11815 $D=1
M59 10 13 VDD VDD P12LL L=1E-07 W=1.2E-06 $X=520 $Y=9005 $D=1
M60 9 32 VDD VDD P12LL L=6E-08 W=5E-07 $X=575 $Y=15760 $D=1
M61 58 VSS VDD VDD P12LL L=2E-07 W=4E-07 $X=585 $Y=2405 $D=1
M62 BLXW[0] 36 VDD VDD P12LL L=6E-08 W=6E-07 $X=610 $Y=16810 $D=1
M63 33 12 57 VDD P12LL L=6E-08 W=4E-07 $X=745 $Y=4300 $D=1
M64 10 CTRCLKW 32 VDD P12LL L=6E-08 W=1.2E-06 $X=790 $Y=10735 $D=1
M65 VDD 32 9 VDD P12LL L=6E-08 W=5E-07 $X=865 $Y=15760 $D=1
M66 VDD 33 10 VDD P12LL L=1E-07 W=1.2E-06 $X=900 $Y=9005 $D=1
M67 BLW[0] 36 BLXW[0] VDD P12LL L=6E-08 W=6E-07 $X=900 $Y=16810 $D=1
M68 17 DATA[0] 58 VDD P12LL L=6E-08 W=4E-07 $X=985 $Y=2405 $D=1
M69 18 35 VDD VDD P12LL L=6E-08 W=5E-07 $X=1155 $Y=15760 $D=1
M70 VDD 36 BLW[0] VDD P12LL L=6E-08 W=6E-07 $X=1190 $Y=16810 $D=1
M71 15 33 VDD VDD P12LL L=1E-07 W=1.2E-06 $X=1270 $Y=9005 $D=1
M72 35 CTRCLKW 15 VDD P12LL L=6E-08 W=1.2E-06 $X=1420 $Y=10735 $D=1
M73 VDD 35 18 VDD P12LL L=6E-08 W=5E-07 $X=1445 $Y=15760 $D=1
M74 VDD 34 34 VDD P12LL L=6E-08 W=4E-07 $X=1480 $Y=4280 $D=1
M75 BLXW[0] 36 VDD VDD P12LL L=6E-08 W=6E-07 $X=1480 $Y=16810 $D=1
M76 VDD VDD DATA[0] VDD P12LL L=6E-08 W=2E-07 $X=1615 $Y=2570 $D=1
M77 VDD 17 15 VDD P12LL L=1E-07 W=1.2E-06 $X=1650 $Y=9005 $D=1
M78 13 17 VDD VDD P12LL L=6E-08 W=4E-07 $X=1760 $Y=4280 $D=1
M79 59 CTRCLKWX 35 VDD P12LL L=6E-08 W=1.2E-07 $X=1760 $Y=11815 $D=1
M80 BLW[0] 36 BLXW[0] VDD P12LL L=6E-08 W=6E-07 $X=1770 $Y=16810 $D=1
M81 VDD 18 59 VDD P12LL L=6E-08 W=1.2E-07 $X=2040 $Y=11815 $D=1
M82 VDD 36 BLW[0] VDD P12LL L=6E-08 W=6E-07 $X=2060 $Y=16810 $D=1
M83 VDD INTCLKX 36 VDD P12LL L=6E-08 W=6E-07 $X=2095 $Y=15725 $D=1
M84 38 INTCLKX VDD VDD P12LL L=6E-08 W=6E-07 $X=2385 $Y=15725 $D=1
M85 BLW[1] 38 VDD VDD P12LL L=6E-08 W=6E-07 $X=2420 $Y=16810 $D=1
M86 60 22 VDD VDD P12LL L=6E-08 W=1.2E-07 $X=2440 $Y=11815 $D=1
M87 BLXW[1] 38 BLW[1] VDD P12LL L=6E-08 W=6E-07 $X=2710 $Y=16810 $D=1
M88 VDD 20 29 VDD P12LL L=6E-08 W=4E-07 $X=2720 $Y=4280 $D=1
M89 39 CTRCLKWX 60 VDD P12LL L=6E-08 W=1.2E-07 $X=2720 $Y=11815 $D=1
M90 24 20 VDD VDD P12LL L=1E-07 W=1.2E-06 $X=2790 $Y=9005 $D=1
M91 DATA[1] VDD VDD VDD P12LL L=6E-08 W=2E-07 $X=2865 $Y=2570 $D=1
M92 40 40 VDD VDD P12LL L=6E-08 W=4E-07 $X=3000 $Y=4280 $D=1
M93 VDD 38 BLXW[1] VDD P12LL L=6E-08 W=6E-07 $X=3000 $Y=16810 $D=1
M94 22 39 VDD VDD P12LL L=6E-08 W=5E-07 $X=3035 $Y=15760 $D=1
M95 24 CTRCLKW 39 VDD P12LL L=6E-08 W=1.2E-06 $X=3060 $Y=10735 $D=1
M96 VDD 41 24 VDD P12LL L=1E-07 W=1.2E-06 $X=3170 $Y=9005 $D=1
M97 BLW[1] 38 VDD VDD P12LL L=6E-08 W=6E-07 $X=3290 $Y=16810 $D=1
M98 VDD 39 22 VDD P12LL L=6E-08 W=5E-07 $X=3325 $Y=15760 $D=1
M99 61 DATA[1] 20 VDD P12LL L=6E-08 W=4E-07 $X=3495 $Y=2405 $D=1
M100 27 41 VDD VDD P12LL L=1E-07 W=1.2E-06 $X=3540 $Y=9005 $D=1
M101 BLXW[1] 38 BLW[1] VDD P12LL L=6E-08 W=6E-07 $X=3580 $Y=16810 $D=1
M102 31 42 VDD VDD P12LL L=6E-08 W=5E-07 $X=3615 $Y=15760 $D=1
M103 42 CTRCLKW 27 VDD P12LL L=6E-08 W=1.2E-06 $X=3690 $Y=10735 $D=1
M104 62 26 41 VDD P12LL L=6E-08 W=4E-07 $X=3735 $Y=4300 $D=1
M105 VDD VSS 61 VDD P12LL L=2E-07 W=4E-07 $X=3755 $Y=2405 $D=1
M106 VDD 38 BLXW[1] VDD P12LL L=6E-08 W=6E-07 $X=3870 $Y=16810 $D=1
M107 VDD 42 31 VDD P12LL L=6E-08 W=5E-07 $X=3905 $Y=15760 $D=1
M108 VDD 29 27 VDD P12LL L=1E-07 W=1.2E-06 $X=3920 $Y=9005 $D=1
M109 63 CTRCLKWX 42 VDD P12LL L=6E-08 W=1.2E-07 $X=4030 $Y=11815 $D=1
M110 VDD VSS 62 VDD P12LL L=2E-07 W=4E-07 $X=4200 $Y=4300 $D=1
M111 VDD 31 63 VDD P12LL L=6E-08 W=1.2E-07 $X=4310 $Y=11815 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: X64Y1D2                                                             *
*******************************************************************************
.SUBCKT qspi_data_info_32_memX64Y1D2 VDD VSS DOUT[1] DOUT[0] BWEN[1] BWEN[0] CTRCLKW CTRCLKWX DIN[1] DIN[0] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] WLA[62] WLA[61] 
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] 
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] 
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] 
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] 
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] 
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] 
+WLA[0] WLB[63] WLB[62] WLB[61] 
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] 
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] 
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] 
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] 
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] 
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] 
+WLB[0] CK1 CK4
XI3 VDD VSS BLA[1] BLA[0] BLXA[1] BLXA[0] DOUT[1] DOUT[0]
+CK1 CK4 qspi_data_info_32_memYMX1R
XI2 VDD VSS BLB[1] BLB[0] BLXB[1] BLXB[0] BWEN[1] BWEN[0] CTRCLKW CTRCLKWX DIN[1] DIN[0] INTCLKX
+qspi_data_info_32_memYMX1W
XI0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0]
+BLXA[1] BLXA[0] BLXB[1] BLXB[0] RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+qspi_data_info_32_memARRAY64X1
.ENDS qspi_data_info_32_memX64Y1D2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TPRF_X64Y1D16                                                       *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTPRF_X64Y1D16 VDD VSS DOUT[15] DOUT[14] DOUT[13] DOUT[12] DOUT[11] 
+DOUT[10] DOUT[9] DOUT[8] DOUT[7] DOUT[6] DOUT[5] DOUT[4] DOUT[3] DOUT[2] DOUT[1] 
+DOUT[0] BWEN[15] BWEN[14] BWEN[13] BWEN[12] BWEN[11] 
+BWEN[10] BWEN[9] BWEN[8] BWEN[7] BWEN[6] BWEN[5] BWEN[4] BWEN[3] BWEN[2] BWEN[1] 
+BWEN[0] CK1 CK4 CTRCLKW CTRCLKWX DIN[15] DIN[14] DIN[13] DIN[12] DIN[11] 
+DIN[10] DIN[9] DIN[8] DIN[7] DIN[6] DIN[5] DIN[4] DIN[3] DIN[2] DIN[1] 
+DIN[0] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1] WLA[63] WLA[62] WLA[61] 
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] 
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] 
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] 
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] 
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] 
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] 
+WLA[0] WLB[63] WLB[62] WLB[61] 
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] 
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] 
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] 
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] 
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] 
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] 
+WLB[0] 
XI2 VDD VSS RWLA[0] RWLA[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+qspi_data_info_32_memTP_EDGECELL64AB
XI1 VDD VSS RWLA[0] RWLA[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+qspi_data_info_32_memTP_EDGECELL64AB
XI0_15 VDD VSS DOUT[15] DOUT[14] BWEN[15] BWEN[14] CTRCLKW CTRCLKWX DIN[15] DIN[14] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_13 VDD VSS DOUT[13] DOUT[12] BWEN[13] BWEN[12] CTRCLKW CTRCLKWX DIN[13] DIN[12] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_11 VDD VSS DOUT[11] DOUT[10] BWEN[11] BWEN[10] CTRCLKW CTRCLKWX DIN[11] DIN[10] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_9 VDD VSS DOUT[9] DOUT[8] BWEN[9] BWEN[8] CTRCLKW CTRCLKWX DIN[9] DIN[8] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_7 VDD VSS DOUT[7] DOUT[6] BWEN[7] BWEN[6] CTRCLKW CTRCLKWX DIN[7] DIN[6] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_5 VDD VSS DOUT[5] DOUT[4] BWEN[5] BWEN[4] CTRCLKW CTRCLKWX DIN[5] DIN[4] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_3 VDD VSS DOUT[3] DOUT[2] BWEN[3] BWEN[2] CTRCLKW CTRCLKWX DIN[3] DIN[2] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_1 VDD VSS DOUT[1] DOUT[0] BWEN[1] BWEN[0] CTRCLKW CTRCLKWX DIN[1] DIN[0] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
.ENDS qspi_data_info_32_memTPRF_X64Y1D16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST                                                        *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST VDD VSS BA BB BXA BXB WLA
*.NOPIN VSS
*.PININFO BA:B BB:B BXA:B BXB:B WLA:I 
MTD0 VSS BCN BC VSS RFNPDHVT W=0.46U L=0.07U M=1
MN2 BXB VSS BCN VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTA1 BXA WLA BCN VSS RFNPGBHVT W=0.12U L=0.09U M=1
MN1 BC VSS BB VSS RFNPGBHVT W=0.12U L=0.09U M=1
MTA0 BC WLA BA VSS RFNPGAHVT W=0.12U L=0.09U M=1
MTD1 BCN BC VSS VSS RFNPDHVT W=0.46U L=0.07U M=1
MTL1 VDD BC BCN VDD RFPLHVT W=0.095U L=0.07U M=1
MTL0 BC BCN VDD VDD RFPLHVT W=0.095U L=0.07U M=1
.ENDS qspi_data_info_32_memTP_BITCELL_ST


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST8A                                                      *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST8A VDD VSS BA0 BA7 BXA0 BXA7 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BA0:B BA7:B BXA0:B BXA7:B DUM_BL:B WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS BA7 DUM_BL BXA7 NET042 WLA[7] qspi_data_info_32_memTP_BITCELL_ST
XI6 VDD VSS NET55 DUM_BL NET54 NET042 WLA[6] qspi_data_info_32_memTP_BITCELL_ST
XI5 VDD VSS NET55 DUM_BL NET54 NET052 WLA[5] qspi_data_info_32_memTP_BITCELL_ST
XI4 VDD VSS NET65 DUM_BL NET64 NET052 WLA[4] qspi_data_info_32_memTP_BITCELL_ST
XI3 VDD VSS NET65 DUM_BL NET64 NET062 WLA[3] qspi_data_info_32_memTP_BITCELL_ST
XI2 VDD VSS NET75 DUM_BL NET74 NET062 WLA[2] qspi_data_info_32_memTP_BITCELL_ST
XI1 VDD VSS NET75 DUM_BL NET74 NET072 WLA[1] qspi_data_info_32_memTP_BITCELL_ST
XI0 VDD VSS BA0 DUM_BL BXA0 NET072 WLA[0] qspi_data_info_32_memTP_BITCELL_ST
.ENDS qspi_data_info_32_memTP_BITCELL_ST8A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BITCELLB2X1                                                          *
*******************************************************************************
.SUBCKT qspi_data_info_32_memBITCELLB2X1 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0]
+WLA[1] WLA[0] WLB[1] WLB[0]
*.NOPIN VSS
*.PININFO BLA[1]:B BLA[0]:B BLB[1]:B BLB[0]:B BLXA[1]:B BLXA[0]:B BLXB[1]:B
*.PININFO BLXB[0]:B WLA[1]:I WLA[0]:I WLB[1]:I WLB[0]:I 
XI0 VDD VSS BLA[1] BLA[0] BLB[1] BLB[0] BLXA[1] BLXA[0] BLXB[1] BLXB[0] WLA[0] WLA[1]
+WLB[0] WLB[1] qspi_data_info_32_memBITCELL2X2
.ENDS qspi_data_info_32_memBITCELLB2X1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST34B                                                     *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST34B VDD VSS DUM_BL RWL[0] RWL[1] WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO DUM_BL:B RWL[0]:I RWL[1]:I WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I
*.PININFO WLA[27]:I WLA[26]:I WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I
*.PININFO WLA[20]:I WLA[19]:I WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I
*.PININFO WLA[13]:I WLA[12]:I WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I
*.PININFO WLA[6]:I WLA[5]:I WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI21 VDD VSS NET035 NET032 qspi_data_info_32_memBLSTRAP_B
XI28 VDD VSS NET056 NET0132 qspi_data_info_32_memBLSTRAP_B
XI26 VDD VSS NET072 DUM_BL NET071 NET064 RWL[1] qspi_data_info_32_memTP_BITCELL_ST
XI27 VDD VSS NET056 DUM_BL NET0132 NET064 RWL[0] qspi_data_info_32_memTP_BITCELL_ST
XI22 VDD VSS NET072 NET051 NET071 NET054 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0] qspi_data_info_32_memTP_BITCELL_ST8A
XI23 VDD VSS NET047 NET051 NET044 NET054 DUM_BL WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] qspi_data_info_32_memTP_BITCELL_ST8A
XI24 VDD VSS NET047 NET039 NET044 NET0130 DUM_BL WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] qspi_data_info_32_memTP_BITCELL_ST8A
XI25 VDD VSS NET035 NET039 NET032 NET0130 DUM_BL WLA[31] WLA[30] WLA[29] WLA[28]
+WLA[27] WLA[26] WLA[25] WLA[24] qspi_data_info_32_memTP_BITCELL_ST8A
.ENDS qspi_data_info_32_memTP_BITCELL_ST34B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST32B                                                     *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST32B VDD VSS DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO DUM_BL:B WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I WLA[26]:I
*.PININFO WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I WLA[19]:I
*.PININFO WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I WLA[12]:I
*.PININFO WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI21 VDD VSS NET45 NET42 qspi_data_info_32_memBLSTRAP_B
XI28 VDD VSS NET66 NET65 qspi_data_info_32_memBLSTRAP_B
XI22 VDD VSS NET66 NET61 NET65 NET64 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] qspi_data_info_32_memTP_BITCELL_ST8A
XI23 VDD VSS NET57 NET61 NET54 NET64 DUM_BL WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] qspi_data_info_32_memTP_BITCELL_ST8A
XI24 VDD VSS NET57 NET49 NET54 NET52 DUM_BL WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] qspi_data_info_32_memTP_BITCELL_ST8A
XI25 VDD VSS NET45 NET49 NET42 NET52 DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] qspi_data_info_32_memTP_BITCELL_ST8A
.ENDS qspi_data_info_32_memTP_BITCELL_ST32B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST8B                                                      *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST8B VDD VSS BXB0 BXB7 DUMBL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BXB0:B BXB7:B DUMBL:B WLA[7]:I WLA[6]:I WLA[5]:I WLA[4]:I WLA[3]:I
*.PININFO WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS NET044 DUMBL NET53 BXB7 WLA[7] qspi_data_info_32_memTP_BITCELL_ST
XI6 VDD VSS NET044 DUMBL NET53 NET045 WLA[6] qspi_data_info_32_memTP_BITCELL_ST
XI5 VDD VSS NET054 DUMBL NET59 NET045 WLA[5] qspi_data_info_32_memTP_BITCELL_ST
XI4 VDD VSS NET054 DUMBL NET59 NET055 WLA[4] qspi_data_info_32_memTP_BITCELL_ST
XI3 VDD VSS NET064 DUMBL NET71 NET055 WLA[3] qspi_data_info_32_memTP_BITCELL_ST
XI2 VDD VSS NET064 DUMBL NET71 NET065 WLA[2] qspi_data_info_32_memTP_BITCELL_ST
XI1 VDD VSS NET074 DUMBL NET83 NET065 WLA[1] qspi_data_info_32_memTP_BITCELL_ST
XI0 VDD VSS NET074 DUMBL NET83 BXB0 WLA[0] qspi_data_info_32_memTP_BITCELL_ST
.ENDS qspi_data_info_32_memTP_BITCELL_ST8B


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST32A                                                     *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST32A VDD VSS DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO DUM_BL:B WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I WLA[26]:I
*.PININFO WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I WLA[19]:I
*.PININFO WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I WLA[12]:I
*.PININFO WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI17 VDD VSS DUM_BL NET47 qspi_data_info_32_memBLSTRAP_A
XI16 VDD VSS DUM_BL NET037 qspi_data_info_32_memBLSTRAP_A
XI0 VDD VSS NET037 NET42 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+qspi_data_info_32_memTP_BITCELL_ST8B
XI1 VDD VSS NET39 NET42 DUM_BL WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] qspi_data_info_32_memTP_BITCELL_ST8B
XI3 VDD VSS NET47 NET34 DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25]
+WLA[24] qspi_data_info_32_memTP_BITCELL_ST8B
XI2 VDD VSS NET39 NET34 DUM_BL WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] qspi_data_info_32_memTP_BITCELL_ST8B
.ENDS qspi_data_info_32_memTP_BITCELL_ST32A


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST8A_TW                                                   *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST8A_TW VDD VSS BA0 BA7 BXA0 BXA7 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4]
+WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BA0:B BA7:B BXA0:B BXA7:B DUM_BL:B WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS BA7 NET043 BXA7 DUM_BL WLA[7] qspi_data_info_32_memTP_BITCELL_ST
XI6 VDD VSS NET55 NET043 NET54 DUM_BL WLA[6] qspi_data_info_32_memTP_BITCELL_ST
XI5 VDD VSS NET55 NET053 NET54 DUM_BL WLA[5] qspi_data_info_32_memTP_BITCELL_ST
XI4 VDD VSS NET65 NET053 NET64 DUM_BL WLA[4] qspi_data_info_32_memTP_BITCELL_ST
XI3 VDD VSS NET65 NET063 NET64 DUM_BL WLA[3] qspi_data_info_32_memTP_BITCELL_ST
XI2 VDD VSS NET75 NET063 NET74 DUM_BL WLA[2] qspi_data_info_32_memTP_BITCELL_ST
XI1 VDD VSS NET75 NET073 NET74 DUM_BL WLA[1] qspi_data_info_32_memTP_BITCELL_ST
XI0 VDD VSS BA0 NET073 BXA0 DUM_BL WLA[0] qspi_data_info_32_memTP_BITCELL_ST
.ENDS qspi_data_info_32_memTP_BITCELL_ST8A_TW


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST32B_TW                                                  *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST32B_TW VDD VSS DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO DUM_BL:B WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I WLA[26]:I
*.PININFO WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I WLA[19]:I
*.PININFO WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I WLA[12]:I
*.PININFO WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI21 VDD VSS NET25 NET22 qspi_data_info_32_memBLSTRAP_B
XI28 VDD VSS NET46 NET45 qspi_data_info_32_memBLSTRAP_B
XI25 VDD VSS NET25 NET29 NET22 NET32 DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] qspi_data_info_32_memTP_BITCELL_ST8A_TW
XI24 VDD VSS NET37 NET29 NET34 NET32 DUM_BL WLA[23] WLA[22] WLA[21] WLA[20] WLA[19]
+WLA[18] WLA[17] WLA[16] qspi_data_info_32_memTP_BITCELL_ST8A_TW
XI22 VDD VSS NET46 NET41 NET45 NET44 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2]
+WLA[1] WLA[0] qspi_data_info_32_memTP_BITCELL_ST8A_TW
XI23 VDD VSS NET37 NET41 NET34 NET44 DUM_BL WLA[15] WLA[14] WLA[13] WLA[12] WLA[11]
+WLA[10] WLA[9] WLA[8] qspi_data_info_32_memTP_BITCELL_ST8A_TW
.ENDS qspi_data_info_32_memTP_BITCELL_ST32B_TW


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST8B_TW                                                   *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST8B_TW VDD VSS BXB0 BXB7 DUMBL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3]
+WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO BXB0:B BXB7:B DUMBL:B WLA[7]:I WLA[6]:I WLA[5]:I WLA[4]:I WLA[3]:I
*.PININFO WLA[2]:I WLA[1]:I WLA[0]:I 
XI7 VDD VSS NET044 BXB7 NET53 DUMBL WLA[7] qspi_data_info_32_memTP_BITCELL_ST
XI6 VDD VSS NET044 NET046 NET53 DUMBL WLA[6] qspi_data_info_32_memTP_BITCELL_ST
XI5 VDD VSS NET054 NET046 NET59 DUMBL WLA[5] qspi_data_info_32_memTP_BITCELL_ST
XI4 VDD VSS NET054 NET056 NET59 DUMBL WLA[4] qspi_data_info_32_memTP_BITCELL_ST
XI3 VDD VSS NET064 NET056 NET71 DUMBL WLA[3] qspi_data_info_32_memTP_BITCELL_ST
XI2 VDD VSS NET064 NET066 NET71 DUMBL WLA[2] qspi_data_info_32_memTP_BITCELL_ST
XI1 VDD VSS NET074 NET066 NET83 DUMBL WLA[1] qspi_data_info_32_memTP_BITCELL_ST
XI0 VDD VSS NET074 BXB0 NET83 DUMBL WLA[0] qspi_data_info_32_memTP_BITCELL_ST
.ENDS qspi_data_info_32_memTP_BITCELL_ST8B_TW


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_BITCELL_ST32A_TW                                                  *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_BITCELL_ST32A_TW VDD VSS DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27]
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8]
+WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
*.NOPIN VSS
*.PININFO DUM_BL:B WLA[31]:I WLA[30]:I WLA[29]:I WLA[28]:I WLA[27]:I WLA[26]:I
*.PININFO WLA[25]:I WLA[24]:I WLA[23]:I WLA[22]:I WLA[21]:I WLA[20]:I WLA[19]:I
*.PININFO WLA[18]:I WLA[17]:I WLA[16]:I WLA[15]:I WLA[14]:I WLA[13]:I WLA[12]:I
*.PININFO WLA[11]:I WLA[10]:I WLA[9]:I WLA[8]:I WLA[7]:I WLA[6]:I WLA[5]:I
*.PININFO WLA[4]:I WLA[3]:I WLA[2]:I WLA[1]:I WLA[0]:I 
XI17 VDD VSS DUM_BL NET033 qspi_data_info_32_memBLSTRAP_B
XI16 VDD VSS DUM_BL NET83 qspi_data_info_32_memBLSTRAP_B
XI3 VDD VSS NET033 NET054 DUM_BL WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] qspi_data_info_32_memTP_BITCELL_ST8B_TW
XI2 VDD VSS NET037 NET054 DUM_BL WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18]
+WLA[17] WLA[16] qspi_data_info_32_memTP_BITCELL_ST8B_TW
XI1 VDD VSS NET037 NET019 DUM_BL WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9]
+WLA[8] qspi_data_info_32_memTP_BITCELL_ST8B_TW
XI0 VDD VSS NET83 NET019 DUM_BL WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+qspi_data_info_32_memTP_BITCELL_ST8B_TW
.ENDS qspi_data_info_32_memTP_BITCELL_ST32A_TW


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_PCAP_EDGE64AB_ST                                                 *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_PCAP_EDGE64AB_ST VDD VSS DUM_BL RWL[0] RWL[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] 
+WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] 
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] 
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] 
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] 
+WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] 
+WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7] 
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
XI3 VDD VSS DUM_BL RWL[0] RWL[1] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] WLA[26]
+WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] WLA[17]
+WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] WLA[8] WLA[7]
+WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] qspi_data_info_32_memTP_BITCELL_ST34B
XI4_1 VDD VSS DUM_BL WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] 
+WLA[54] WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] 
+WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] 
+WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] qspi_data_info_32_memTP_BITCELL_ST32A_TW
.ENDS qspi_data_info_32_memTP_PCAP_EDGE64AB_ST


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TPRF_X64Y1D16_ST                                                    *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTPRF_X64Y1D16_ST VDD VSS DOUT[15] DOUT[14] DOUT[13] DOUT[12] DOUT[11] 
+DOUT[10] DOUT[9] DOUT[8] DOUT[7] DOUT[6] DOUT[5] DOUT[4] DOUT[3] DOUT[2] DOUT[1] 
+DOUT[0] BWEN[15] BWEN[14] BWEN[13] BWEN[12] BWEN[11] 
+BWEN[10] BWEN[9] BWEN[8] BWEN[7] BWEN[6] BWEN[5] BWEN[4] BWEN[3] BWEN[2] BWEN[1] 
+BWEN[0] CK1 CK4 CTRCLKW CTRCLKWX DBLA DIN[15] DIN[14] DIN[13] DIN[12] DIN[11] 
+DIN[10] DIN[9] DIN[8] DIN[7] DIN[6] DIN[5] DIN[4] DIN[3] DIN[2] DIN[1] 
+DIN[0] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1] WLA[63] WLA[62] WLA[61] 
+WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] 
+WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] 
+WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] 
+WLA[30] WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] 
+WLA[20] WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] 
+WLA[10] WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] 
+WLA[0] WLB[63] WLB[62] WLB[61] 
+WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] 
+WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] 
+WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] 
+WLB[30] WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] 
+WLB[20] WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] 
+WLB[10] WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] 
+WLB[0] 
XI2 VDD VSS RWLA[0] RWLA[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+qspi_data_info_32_memTP_EDGECELL64AB
XI1 VDD VSS DBLA RWLA[0] RWLA[1] WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+qspi_data_info_32_memTP_PCAP_EDGE64AB_ST
XI0_15 VDD VSS DOUT[15] DOUT[14] BWEN[15] BWEN[14] CTRCLKW CTRCLKWX DIN[15] DIN[14] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_13 VDD VSS DOUT[13] DOUT[12] BWEN[13] BWEN[12] CTRCLKW CTRCLKWX DIN[13] DIN[12] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_11 VDD VSS DOUT[11] DOUT[10] BWEN[11] BWEN[10] CTRCLKW CTRCLKWX DIN[11] DIN[10] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_9 VDD VSS DOUT[9] DOUT[8] BWEN[9] BWEN[8] CTRCLKW CTRCLKWX DIN[9] DIN[8] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_7 VDD VSS DOUT[7] DOUT[6] BWEN[7] BWEN[6] CTRCLKW CTRCLKWX DIN[7] DIN[6] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_5 VDD VSS DOUT[5] DOUT[4] BWEN[5] BWEN[4] CTRCLKW CTRCLKWX DIN[5] DIN[4] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_3 VDD VSS DOUT[3] DOUT[2] BWEN[3] BWEN[2] CTRCLKW CTRCLKWX DIN[3] DIN[2] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
XI0_1 VDD VSS DOUT[1] DOUT[0] BWEN[1] BWEN[0] CTRCLKW CTRCLKWX DIN[1] DIN[0] INTCLKX RWLA[0] RWLA[1] RWLB[0] RWLB[1]
+WLA[63] 
+WLA[62] WLA[61] WLA[60] WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] 
+WLA[53] WLA[52] WLA[51] WLA[50] WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] 
+WLA[44] WLA[43] WLA[42] WLA[41] WLA[40] WLA[39] WLA[38] WLA[37] WLA[36] 
+WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30] WLA[29] WLA[28] WLA[27] 
+WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20] WLA[19] WLA[18] 
+WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10] WLA[9] 
+WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0] 
+WLB[63] 
+WLB[62] WLB[61] WLB[60] WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] 
+WLB[53] WLB[52] WLB[51] WLB[50] WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] 
+WLB[44] WLB[43] WLB[42] WLB[41] WLB[40] WLB[39] WLB[38] WLB[37] WLB[36] 
+WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30] WLB[29] WLB[28] WLB[27] 
+WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20] WLB[19] WLB[18] 
+WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10] WLB[9] 
+WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0] 
+CK1 CK4 qspi_data_info_32_memX64Y1D2
.ENDS qspi_data_info_32_memTPRF_X64Y1D16_ST


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: ESDA5W                                                               *
*******************************************************************************
.SUBCKT qspi_data_info_32_memESDA5W VDD VSS A[5] A[4] A[3] A[2] A[1] A[0] 
+CEN CLK
MN5 A[5] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP5 VDD VDD A[5] VDD P12LL W=0.2U L=0.06U M=1
MN4 A[4] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP4 VDD VDD A[4] VDD P12LL W=0.2U L=0.06U M=1
MN3 A[3] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP3 VDD VDD A[3] VDD P12LL W=0.2U L=0.06U M=1
MN2 A[2] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP2 VDD VDD A[2] VDD P12LL W=0.2U L=0.06U M=1
MN1 A[1] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP1 VDD VDD A[1] VDD P12LL W=0.2U L=0.06U M=1
MN0 A[0] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP0 VDD VDD A[0] VDD P12LL W=0.2U L=0.06U M=1
MN123 CEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP123 VDD VDD CEN VDD P12LL W=0.2U L=0.06U M=1
MN120 CLK VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP120 VDD VDD CLK VDD P12LL W=0.2U L=0.06U M=1
.ENDS qspi_data_info_32_memESDA5W


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: ESDA5R                                                               *
*******************************************************************************
.SUBCKT qspi_data_info_32_memESDA5R VDD VSS A[5] A[4] A[3] A[2] A[1] A[0] 
+CEN CLK RDE 
MN5 A[5] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP5 VDD VDD A[5] VDD P12LL W=0.2U L=0.06U M=1
MN4 A[4] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP4 VDD VDD A[4] VDD P12LL W=0.2U L=0.06U M=1
MN3 A[3] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP3 VDD VDD A[3] VDD P12LL W=0.2U L=0.06U M=1
MN2 A[2] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP2 VDD VDD A[2] VDD P12LL W=0.2U L=0.06U M=1
MN1 A[1] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP1 VDD VDD A[1] VDD P12LL W=0.2U L=0.06U M=1
MN0 A[0] VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP0 VDD VDD A[0] VDD P12LL W=0.2U L=0.06U M=1
MN120 CLK VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP120 VDD VDD CLK VDD P12LL W=0.2U L=0.06U M=1
MN127 RDE VSS VSS VSS N12LL W=0.4U L=0.06U M=1
MP127 VDD VDD RDE VDD P12LL W=0.4U L=0.06U M=1
MN123 CEN VSS VSS VSS N12LL W=0.2U L=0.06U M=1
MP123 VDD VDD CEN VDD P12LL W=0.2U L=0.06U M=1
.ENDS qspi_data_info_32_memESDA5R


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: OPDEC                                                                *
*******************************************************************************
.SUBCKT qspi_data_info_32_memOPDEC VDD VSS S[5] S[4] S[3] S[2] S[1] S[0] OP[2] OP[1] OP[0]

M0 VSS OP[0] 21 VSS N12LL L=6E-08 W=4E-07 $X=2670 $Y=4295 $D=0
M1 23 21 VSS VSS N12LL L=6E-08 W=4E-07 $X=2960 $Y=4295 $D=0
M2 VSS OP[1] 26 VSS N12LL L=6E-08 W=4E-07 $X=3665 $Y=4295 $D=0
M3 25 26 VSS VSS N12LL L=6E-08 W=4E-07 $X=3955 $Y=4295 $D=0
M4 37 21 S[0] VSS N12LL L=6E-08 W=4E-07 $X=4880 $Y=4310 $D=0
M5 38 36 37 VSS N12LL L=6E-08 W=4E-07 $X=5170 $Y=4310 $D=0
M6 VSS 26 38 VSS N12LL L=6E-08 W=4E-07 $X=5460 $Y=4310 $D=0
M7 39 26 VSS VSS N12LL L=6E-08 W=4E-07 $X=5755 $Y=4310 $D=0
M8 S[1] 36 39 VSS N12LL L=6E-08 W=4E-07 $X=6045 $Y=4310 $D=0
M9 40 36 S[2] VSS N12LL L=6E-08 W=4E-07 $X=6675 $Y=4310 $D=0
M10 VSS 31 40 VSS N12LL L=6E-08 W=4E-07 $X=6965 $Y=4310 $D=0
M11 41 23 VSS VSS N12LL L=6E-08 W=4E-07 $X=7265 $Y=4310 $D=0
M12 31 25 41 VSS N12LL L=6E-08 W=4E-07 $X=7555 $Y=4310 $D=0
M13 32 25 VSS VSS N12LL L=6E-08 W=4E-07 $X=8185 $Y=4310 $D=0
M14 VSS 23 32 VSS N12LL L=6E-08 W=4E-07 $X=8475 $Y=4310 $D=0
M15 S[4] 32 VSS VSS N12LL L=6E-08 W=4E-07 $X=8775 $Y=4310 $D=0
M16 VSS 36 S[4] VSS N12LL L=6E-08 W=4E-07 $X=9065 $Y=4310 $D=0
M17 S[5] 26 VSS VSS N12LL L=6E-08 W=4E-07 $X=9695 $Y=4310 $D=0
M18 VSS 36 S[5] VSS N12LL L=6E-08 W=4E-07 $X=9985 $Y=4310 $D=0
M19 VSS 36 S[3] VSS N12LL L=6E-08 W=4E-07 $X=10670 $Y=4295 $D=0
M20 36 OP[2] VSS VSS N12LL L=6E-08 W=4E-07 $X=10960 $Y=4295 $D=0
M21 VDD OP[0] 21 VDD P12LL L=6E-08 W=4E-07 $X=2670 $Y=5405 $D=1
M22 23 21 VDD VDD P12LL L=6E-08 W=4E-07 $X=2960 $Y=5405 $D=1
M23 VDD OP[1] 26 VDD P12LL L=6E-08 W=4E-07 $X=3665 $Y=5405 $D=1
M24 25 26 VDD VDD P12LL L=6E-08 W=4E-07 $X=3955 $Y=5405 $D=1
M25 VDD 21 S[0] VDD P12LL L=6E-08 W=4E-07 $X=4880 $Y=5420 $D=1
M26 S[0] 36 VDD VDD P12LL L=6E-08 W=4E-07 $X=5170 $Y=5420 $D=1
M27 VDD 26 S[0] VDD P12LL L=6E-08 W=4E-07 $X=5460 $Y=5420 $D=1
M28 S[1] 26 VDD VDD P12LL L=6E-08 W=4E-07 $X=5755 $Y=5420 $D=1
M29 VDD 36 S[1] VDD P12LL L=6E-08 W=4E-07 $X=6045 $Y=5420 $D=1
M30 S[2] 36 VDD VDD P12LL L=6E-08 W=4E-07 $X=6675 $Y=5420 $D=1
M31 VDD 31 S[2] VDD P12LL L=6E-08 W=4E-07 $X=6965 $Y=5420 $D=1
M32 31 23 VDD VDD P12LL L=6E-08 W=4E-07 $X=7265 $Y=5420 $D=1
M33 VDD 25 31 VDD P12LL L=6E-08 W=4E-07 $X=7555 $Y=5420 $D=1
M34 42 25 32 VDD P12LL L=6E-08 W=4E-07 $X=8185 $Y=5420 $D=1
M35 VDD 23 42 VDD P12LL L=6E-08 W=4E-07 $X=8475 $Y=5420 $D=1
M36 43 32 VDD VDD P12LL L=6E-08 W=4E-07 $X=8775 $Y=5420 $D=1
M37 S[4] 36 43 VDD P12LL L=6E-08 W=4E-07 $X=9065 $Y=5420 $D=1
M38 44 26 S[5] VDD P12LL L=6E-08 W=4E-07 $X=9695 $Y=5420 $D=1
M39 VDD 36 44 VDD P12LL L=6E-08 W=4E-07 $X=9985 $Y=5420 $D=1
M40 VDD 36 S[3] VDD P12LL L=6E-08 W=4E-07 $X=10670 $Y=5425 $D=1
M41 36 OP[2] VDD VDD P12LL L=6E-08 W=4E-07 $X=10960 $Y=5425 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDEC                                                                 *
*******************************************************************************
.SUBCKT qspi_data_info_32_memXDEC VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] FCK[7] FCK[6]
+FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA PXB PXC

M0 25 26 VSS VSS N12LL L=6E-08 W=5.05E-07 $X=2425 $Y=2195 $D=0
M1 VSS 26 25 VSS N12LL L=6E-08 W=5.05E-07 $X=2425 $Y=2485 $D=0
M2 26 23 VSS VSS N12LL L=6E-08 W=5.05E-07 $X=2425 $Y=2775 $D=0
M3 VSS 23 26 VSS N12LL L=6E-08 W=5.05E-07 $X=2425 $Y=3065 $D=0
M4 59 PXC 23 VSS N12LL L=6E-08 W=8.0E-07 $X=2425 $Y=3725 $D=0
M5 60 PXB 59 VSS N12LL L=6E-08 W=8.0E-07 $X=2425 $Y=4015 $D=0
M6 VSS PXA 60 VSS N12LL L=6E-08 W=8.0E-07 $X=2425 $Y=4305 $D=0
M7 FCK[1] 26 28 VSS N12LL L=6E-08 W=7E-07 $X=9360 $Y=1415 $D=0
M8 30 26 FCK[3] VSS N12LL L=6E-08 W=7E-07 $X=9360 $Y=2430 $D=0
M9 FCK[5] 26 32 VSS N12LL L=6E-08 W=7E-07 $X=9360 $Y=3735 $D=0
M10 FCK[7] 26 34 VSS N12LL L=6E-08 W=7E-07 $X=9360 $Y=4725 $D=0
M11 27 26 FCK[0] VSS N12LL L=6E-08 W=7E-07 $X=10285 $Y=910 $D=0
M12 29 26 FCK[2] VSS N12LL L=6E-08 W=7E-07 $X=10285 $Y=1920 $D=0
M13 31 26 FCK[4] VSS N12LL L=6E-08 W=7E-07 $X=10285 $Y=2935 $D=0
M14 FCK[6] 26 33 VSS N12LL L=6E-08 W=7E-07 $X=10285 $Y=4225 $D=0
M15 35 27 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=900 $D=0
M16 VSS 27 35 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=1160 $D=0
M17 36 28 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=1410 $D=0
M18 VSS 28 36 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=1670 $D=0
M19 37 29 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=1920 $D=0
M20 VSS 29 37 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=2180 $D=0
M21 38 30 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=2430 $D=0
M22 VSS 30 38 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=2690 $D=0
M23 39 31 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=2940 $D=0
M24 VSS 31 39 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=3200 $D=0
M25 40 32 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=3450 $D=0
M26 VSS 32 40 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=3710 $D=0
M27 41 33 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=3960 $D=0
M28 VSS 33 41 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=4220 $D=0
M29 42 34 VSS VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=4470 $D=0
M30 VSS 34 42 VSS N12LL L=6E-08 W=5E-07 $X=11625 $Y=4730 $D=0
M31 WL[0] 43 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=900 $D=0
M32 VSS 43 WL[0] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=1160 $D=0
M33 WL[1] 44 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=1410 $D=0
M34 VSS 44 WL[1] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=1670 $D=0
M35 WL[2] 45 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=1920 $D=0
M36 VSS 45 WL[2] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=2180 $D=0
M37 WL[3] 46 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=2430 $D=0
M38 VSS 46 WL[3] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=2690 $D=0
M39 WL[4] 47 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=2940 $D=0
M40 VSS 47 WL[4] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=3200 $D=0
M41 WL[5] 48 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=3450 $D=0
M42 VSS 48 WL[5] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=3710 $D=0
M43 WL[6] 49 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=3960 $D=0
M44 VSS 49 WL[6] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=4220 $D=0
M45 WL[7] 50 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=4470 $D=0
M46 VSS 50 WL[7] VSS N12LL L=6E-08 W=2.5E-06 $X=19190 $Y=4730 $D=0
M47 43 35 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=900 $D=6
M48 VSS 35 43 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=1160 $D=6
M49 44 36 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=1410 $D=6
M50 VSS 36 44 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=1670 $D=6
M51 45 37 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=1920 $D=6
M52 VSS 37 45 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=2180 $D=6
M53 46 38 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=2430 $D=6
M54 VSS 38 46 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=2690 $D=6
M55 47 39 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=2940 $D=6
M56 VSS 39 47 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=3200 $D=6
M57 48 40 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=3450 $D=6
M58 VSS 40 48 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=3710 $D=6
M59 49 41 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=3960 $D=6
M60 VSS 41 49 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=4220 $D=6
M61 50 42 VSS VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=4470 $D=6
M62 VSS 42 50 VSS NHVT12LL L=6E-08 W=1.25E-06 $X=17395 $Y=4730 $D=6
M63 WL[0] 43 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=900 $D=7
M64 VDD 43 WL[0] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=1160 $D=7
M65 WL[1] 44 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=1410 $D=7
M66 VDD 44 WL[1] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=1670 $D=7
M67 WL[2] 45 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=1920 $D=7
M68 VDD 45 WL[2] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=2180 $D=7
M69 WL[3] 46 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=2430 $D=7
M70 VDD 46 WL[3] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=2690 $D=7
M71 WL[4] 47 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=2940 $D=7
M72 VDD 47 WL[4] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=3200 $D=7
M73 WL[5] 48 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=3450 $D=7
M74 VDD 48 WL[5] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=3710 $D=7
M75 WL[6] 49 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=3960 $D=7
M76 VDD 49 WL[6] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=4220 $D=7
M77 WL[7] 50 VDD VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=4470 $D=7
M78 VDD 50 WL[7] VDD PHVT12LL L=6E-08 W=5E-06 $X=22090 $Y=4730 $D=7
M79 25 26 VDD VDD P12LL L=6E-08 W=5E-07 $X=3930 $Y=2195 $D=1
M80 VDD 26 25 VDD P12LL L=6E-08 W=5E-07 $X=3930 $Y=2485 $D=1
M81 26 23 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=3930 $Y=2775 $D=1
M82 VDD 23 26 VDD P12LL L=6E-08 W=7.5E-07 $X=3930 $Y=3065 $D=1
M83 VDD PXC 23 VDD P12LL L=6E-08 W=5E-07 $X=3930 $Y=3725 $D=1
M84 23 PXB VDD VDD P12LL L=6E-08 W=5E-07 $X=3930 $Y=4015 $D=1
M85 VDD PXA 23 VDD P12LL L=6E-08 W=5E-07 $X=3930 $Y=4305 $D=1
M86 27 26 VDD VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=910 $D=1
M87 VDD 26 28 VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=1490 $D=1
M88 29 26 VDD VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=1770 $D=1
M89 VDD 26 30 VDD P12LL L=6E-08 W=5.15E-07 $X=6070 $Y=2700 $D=1
M90 31 26 VDD VDD P12LL L=6E-08 W=5.15E-07 $X=6070 $Y=2970 $D=1
M91 VDD 26 32 VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=3820 $D=1
M92 33 26 VDD VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=4100 $D=1
M93 VDD 26 34 VDD P12LL L=6E-08 W=5E-07 $X=6070 $Y=4725 $D=1
M94 FCK[1] 25 28 VDD P12LL L=6E-08 W=4E-07 $X=7195 $Y=1415 $D=1
M95 30 25 FCK[3] VDD P12LL L=6E-08 W=4E-07 $X=7195 $Y=2585 $D=1
M96 FCK[5] 25 32 VDD P12LL L=6E-08 W=4E-07 $X=7195 $Y=3730 $D=1
M97 FCK[7] 25 34 VDD P12LL L=6E-08 W=4E-07 $X=7195 $Y=4725 $D=1
M98 27 25 FCK[0] VDD P12LL L=6E-08 W=4E-07 $X=8015 $Y=910 $D=1
M99 29 25 FCK[2] VDD P12LL L=6E-08 W=4E-07 $X=8015 $Y=1920 $D=1
M100 FCK[6] 25 33 VDD P12LL L=6E-08 W=4E-07 $X=8015 $Y=4225 $D=1
M101 31 25 FCK[4] VDD P12LL L=6E-08 W=4E-07 $X=8055 $Y=2950 $D=1
M102 35 27 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=900 $D=1
M103 VDD 27 35 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=1160 $D=1
M104 36 28 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=1410 $D=1
M105 VDD 28 36 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=1670 $D=1
M106 37 29 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=1920 $D=1
M107 VDD 29 37 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=2180 $D=1
M108 38 30 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=2430 $D=1
M109 VDD 30 38 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=2690 $D=1
M110 39 31 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=2940 $D=1
M111 VDD 31 39 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=3200 $D=1
M112 40 32 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=3450 $D=1
M113 VDD 32 40 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=3710 $D=1
M114 41 33 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=3960 $D=1
M115 VDD 33 41 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=4220 $D=1
M116 42 34 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=4470 $D=1
M117 VDD 34 42 VDD P12LL L=6E-08 W=1.25E-06 $X=12625 $Y=4730 $D=1
M118 43 35 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=900 $D=1
M119 VDD 35 43 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=1160 $D=1
M120 44 36 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=1410 $D=1
M121 VDD 36 44 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=1670 $D=1
M122 45 37 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=1920 $D=1
M123 VDD 37 45 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=2180 $D=1
M124 46 38 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=2430 $D=1
M125 VDD 38 46 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=2690 $D=1
M126 47 39 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=2940 $D=1
M127 VDD 39 47 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=3200 $D=1
M128 48 40 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=3450 $D=1
M129 VDD 40 48 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=3710 $D=1
M130 49 41 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=3960 $D=1
M131 VDD 41 49 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=4220 $D=1
M132 50 42 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=4470 $D=1
M133 VDD 42 50 VDD P12LL L=6E-08 W=2.5E-06 $X=14395 $Y=4730 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDEC8                                                               *
*******************************************************************************
.SUBCKT qspi_data_info_32_memXDEC8 VDD VSS WL[63] 
+WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] 
+WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] 
+WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] 
+WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] 
+WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] 
+WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] 
+WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0]
+PXA[3] PXA[2] PXA[1] PXA[0] PXB[1] PXB[0] PXC[0]
XI86_7 VDD VSS WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[3] PXB[1] PXC[0] qspi_data_info_32_memXDEC
XI86_6 VDD VSS WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[2] PXB[1] PXC[0] qspi_data_info_32_memXDEC
XI86_5 VDD VSS WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[1] PXB[1] PXC[0] qspi_data_info_32_memXDEC
XI86_4 VDD VSS WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[0] PXB[1] PXC[0] qspi_data_info_32_memXDEC
XI86_3 VDD VSS WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[3] PXB[0] PXC[0] qspi_data_info_32_memXDEC
XI86_2 VDD VSS WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[2] PXB[0] PXC[0] qspi_data_info_32_memXDEC
XI86_1 VDD VSS WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[1] PXB[0] PXC[0] qspi_data_info_32_memXDEC
XI86_0 VDD VSS WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] 
+FCK[7] FCK[6] FCK[5] FCK[4] FCK[3] FCK[2] FCK[1] FCK[0] PXA[0] PXB[0] PXC[0] qspi_data_info_32_memXDEC
.ENDS qspi_data_info_32_memXDEC8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_CLKW                                                              *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_CLKW VDD VSS ACTRCLK ACTRCLKX DCTRCLK DCTRCLKX INTCLKX CEN CLK
* SPICE NETLIST

M0 35 34 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=405 $Y=9475 $D=0
M1 VSS 34 35 VSS N12LL L=6E-08 W=1.25E-06 $X=695 $Y=9475 $D=0
M2 34 21 VSS VSS N12LL L=6E-08 W=8E-07 $X=985 $Y=9925 $D=0
M3 36 CLK VSS VSS N12LL L=6E-08 W=4E-07 $X=1715 $Y=3545 $D=0
M4 21 37 VSS VSS N12LL L=6E-08 W=6.05E-07 $X=1765 $Y=9995 $D=0
M5 VSS 37 21 VSS N12LL L=6E-08 W=6.05E-07 $X=2055 $Y=9995 $D=0
M6 37 40 VSS VSS N12LL L=6E-08 W=1E-06 $X=2355 $Y=9600 $D=0
M7 85 36 VSS VSS N12LL L=6E-08 W=1E-06 $X=2365 $Y=3540 $D=0
M8 39 CEN 85 VSS N12LL L=6E-08 W=1E-06 $X=2605 $Y=3540 $D=0
M9 VSS 40 37 VSS N12LL L=6E-08 W=1E-06 $X=2640 $Y=9600 $D=0
M10 VSS 52 39 VSS N12LL L=6E-07 W=1.2E-07 $X=3275 $Y=3830 $D=0
M11 86 VDD 40 VSS N12LL L=4E-07 W=8E-07 $X=3355 $Y=9665 $D=0
M12 VSS 39 52 VSS N12LL L=6E-08 W=4E-07 $X=3920 $Y=3615 $D=0
M13 VSS 41 86 VSS N12LL L=6E-08 W=8E-07 $X=3955 $Y=9665 $D=0
M14 42 52 VSS VSS N12LL L=6E-08 W=5E-07 $X=4210 $Y=3615 $D=0
M15 51 CLK 22 VSS N12LL L=6E-08 W=4E-06 $X=4280 $Y=4970 $D=0
M16 41 43 VSS VSS N12LL L=2E-07 W=4E-07 $X=4305 $Y=10065 $D=0
M17 VSS CLK 42 VSS N12LL L=6E-08 W=5E-07 $X=4500 $Y=3615 $D=0
M18 22 CLK 51 VSS N12LL L=6E-08 W=4E-06 $X=4570 $Y=4970 $D=0
M19 51 CLK 22 VSS N12LL L=6E-08 W=4E-06 $X=4860 $Y=4970 $D=0
M20 22 CLK 51 VSS N12LL L=6E-08 W=4E-06 $X=5150 $Y=4970 $D=0
M21 VSS 42 44 VSS N12LL L=6E-08 W=5E-07 $X=5190 $Y=3495 $D=0
M22 VSS 45 43 VSS N12LL L=2E-07 W=4E-07 $X=5405 $Y=10220 $D=0
M23 51 CLK 22 VSS N12LL L=6E-08 W=4E-06 $X=5440 $Y=4970 $D=0
M24 46 44 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5540 $Y=3495 $D=0
M25 VSS 44 46 VSS N12LL L=6E-08 W=7.5E-07 $X=5830 $Y=3495 $D=0
M26 45 47 VSS VSS N12LL L=2E-07 W=4E-07 $X=5935 $Y=10220 $D=0
M27 51 46 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=6100 $Y=6125 $D=0
M28 VSS 46 51 VSS N12LL L=6E-08 W=2.5E-06 $X=6390 $Y=6125 $D=0
M29 51 46 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=6680 $Y=6125 $D=0
M30 VSS 50 47 VSS N12LL L=2E-07 W=4E-07 $X=6850 $Y=10220 $D=0
M31 VSS 46 51 VSS N12LL L=6E-08 W=2.5E-06 $X=6970 $Y=6125 $D=0
M32 51 46 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=7260 $Y=6125 $D=0
M33 50 22 VSS VSS N12LL L=6E-08 W=7E-07 $X=7340 $Y=9920 $D=0
M34 VSS 46 51 VSS N12LL L=6E-08 W=2.5E-06 $X=7550 $Y=6125 $D=0
M35 51 46 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=7840 $Y=6125 $D=0
M36 VSS 53 25 VSS N12LL L=2E-07 W=4E-07 $X=7895 $Y=3465 $D=0
M37 VSS 46 51 VSS N12LL L=6E-08 W=2.5E-06 $X=8130 $Y=6125 $D=0
M38 53 VSS VSS VSS N12LL L=2E-07 W=4E-07 $X=8395 $Y=3465 $D=0
M39 54 25 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=8420 $Y=6125 $D=0
M40 VSS 58 54 VSS N12LL L=6E-08 W=2.5E-06 $X=8710 $Y=6125 $D=0
M41 VSS 58 53 VSS N12LL L=2E-07 W=4E-07 $X=8905 $Y=3465 $D=0
M42 ACTRCLK 54 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=9000 $Y=6125 $D=0
M43 VSS 54 ACTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=9290 $Y=6125 $D=0
M44 DCTRCLK 54 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=9580 $Y=6125 $D=0
M45 VSS 54 DCTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=9870 $Y=6125 $D=0
M46 VSS 58 22 VSS N12LL L=1E-06 W=1.2E-07 $X=10120 $Y=4325 $D=0
M47 ACTRCLKX ACTRCLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=10160 $Y=6125 $D=0
M48 VSS ACTRCLK ACTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=10450 $Y=6125 $D=0
M49 DCTRCLKX 30 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=10740 $Y=6125 $D=0
M50 VSS 30 DCTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=11030 $Y=6125 $D=0
M51 30 54 VSS VSS N12LL L=6E-08 W=3E-06 $X=11310 $Y=5625 $D=0
M52 58 22 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=11900 $Y=6125 $D=0
M53 VSS 22 58 VSS N12LL L=6E-08 W=2.5E-06 $X=12190 $Y=6125 $D=0
M54 58 22 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=12480 $Y=6125 $D=0
M55 VSS 22 58 VSS N12LL L=6E-08 W=2.5E-06 $X=12770 $Y=6125 $D=0
M56 INTCLKX 58 VSS VSS N12LL L=6E-08 W=5E-06 $X=13640 $Y=3625 $D=0
M57 VSS 57 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=13930 $Y=3625 $D=0
M58 INTCLKX 57 VSS VSS N12LL L=6E-08 W=5E-06 $X=14220 $Y=3625 $D=0
M59 VSS 58 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=14510 $Y=3625 $D=0
M60 INTCLKX 58 VSS VSS N12LL L=6E-08 W=5E-06 $X=14800 $Y=3625 $D=0
M61 VSS 57 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=15090 $Y=3625 $D=0
M62 INTCLKX 57 VSS VSS N12LL L=6E-08 W=5E-06 $X=15380 $Y=3625 $D=0
M63 VSS 58 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=15670 $Y=3625 $D=0
M64 57 59 VSS VSS N12LL L=6E-08 W=7E-07 $X=15990 $Y=3625 $D=0
M65 VSS 59 57 VSS N12LL L=6E-08 W=7E-07 $X=16280 $Y=3625 $D=0
M66 59 58 VSS VSS N12LL L=6E-08 W=4E-07 $X=16570 $Y=3625 $D=0
M67 35 34 VDD VDD P12LL L=6E-08 W=1.24E-06 $X=405 $Y=11385 $D=2
M68 VDD 34 35 VDD P12LL L=6E-08 W=1.24E-06 $X=695 $Y=11385 $D=2
M69 34 21 VDD VDD P12LL L=6E-08 W=8E-07 $X=985 $Y=11385 $D=2
M70 36 CLK VDD VDD P12LL L=6E-08 W=4E-07 $X=1715 $Y=2250 $D=2
M71 21 37 VDD VDD P12LL L=6E-08 W=1.2E-06 $X=1765 $Y=11385 $D=2
M72 VDD 37 21 VDD P12LL L=6E-08 W=1.2E-06 $X=2055 $Y=11385 $D=2
M73 37 40 VDD VDD P12LL L=6E-08 W=2E-06 $X=2355 $Y=11385 $D=2
M74 91 CLK VDD VDD P12LL L=6E-08 W=1E-06 $X=2365 $Y=1670 $D=2
M75 39 CEN 91 VDD P12LL L=6E-08 W=1E-06 $X=2605 $Y=1670 $D=2
M76 VDD 40 37 VDD P12LL L=6E-08 W=2E-06 $X=2640 $Y=11385 $D=2
M77 VDD 52 39 VDD P12LL L=3E-07 W=1.2E-07 $X=2975 $Y=2435 $D=2
M78 92 VSS 40 VDD P12LL L=4E-07 W=1.2E-06 $X=3355 $Y=11355 $D=2
M79 21 50 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=3845 $Y=13320 $D=2
M80 VDD 39 52 VDD P12LL L=6E-08 W=8E-07 $X=3920 $Y=1870 $D=2
M81 VDD 41 92 VDD P12LL L=6E-08 W=1.2E-06 $X=3955 $Y=11355 $D=2
M82 VDD 50 21 VDD P12LL L=6E-08 W=1.25E-06 $X=4135 $Y=13320 $D=2
M83 93 52 VDD VDD P12LL L=6E-08 W=1E-06 $X=4210 $Y=1670 $D=2
M84 41 43 VDD VDD P12LL L=2E-07 W=6E-07 $X=4305 $Y=11355 $D=2
M85 22 35 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=4425 $Y=13320 $D=2
M86 42 CLK 93 VDD P12LL L=6E-08 W=1E-06 $X=4500 $Y=1670 $D=2
M87 VDD 35 22 VDD P12LL L=6E-08 W=1.25E-06 $X=4715 $Y=13320 $D=2
M88 22 35 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5005 $Y=13320 $D=2
M89 VDD 42 44 VDD P12LL L=6E-08 W=1E-06 $X=5190 $Y=1800 $D=2
M90 VDD 35 22 VDD P12LL L=6E-08 W=1.25E-06 $X=5295 $Y=13320 $D=2
M91 VDD 45 43 VDD P12LL L=2E-07 W=6E-07 $X=5405 $Y=11385 $D=2
M92 46 44 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=5540 $Y=1300 $D=2
M93 22 35 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5585 $Y=13320 $D=2
M94 VDD 44 46 VDD P12LL L=6E-08 W=1.5E-06 $X=5830 $Y=1300 $D=2
M95 VDD 35 22 VDD P12LL L=6E-08 W=1.25E-06 $X=5875 $Y=13320 $D=2
M96 45 47 VDD VDD P12LL L=2E-07 W=6E-07 $X=5935 $Y=11385 $D=2
M97 22 35 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=6165 $Y=13320 $D=2
M98 VDD 35 22 VDD P12LL L=6E-08 W=1.25E-06 $X=6455 $Y=13320 $D=2
M99 VDD 50 47 VDD P12LL L=2E-07 W=6E-07 $X=6850 $Y=11385 $D=2
M100 50 22 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=7340 $Y=11385 $D=2
M101 VDD 53 25 VDD P12LL L=2E-07 W=4E-07 $X=7895 $Y=2040 $D=2
M102 97 VSS VDD VDD P12LL L=2E-07 W=8E-07 $X=8395 $Y=2040 $D=2
M103 96 25 54 VDD P12LL L=6E-08 W=2.5E-06 $X=8420 $Y=9420 $D=2
M104 VDD 58 96 VDD P12LL L=6E-08 W=2.5E-06 $X=8660 $Y=9420 $D=2
M105 53 58 97 VDD P12LL L=2E-07 W=8E-07 $X=8905 $Y=2040 $D=2
M106 ACTRCLK 54 VDD VDD P12LL L=6E-08 W=5E-06 $X=9000 $Y=9420 $D=2
M107 VDD 54 ACTRCLK VDD P12LL L=6E-08 W=5E-06 $X=9290 $Y=9420 $D=2
M108 DCTRCLK 54 VDD VDD P12LL L=6E-08 W=5E-06 $X=9580 $Y=9420 $D=2
M109 VDD 54 DCTRCLK VDD P12LL L=6E-08 W=5E-06 $X=9870 $Y=9420 $D=2
M110 ACTRCLKX ACTRCLK VDD VDD P12LL L=6E-08 W=5E-06 $X=10160 $Y=9420 $D=2
M111 22 58 VDD VDD P12LL L=2E-07 W=1.2E-07 $X=10215 $Y=2370 $D=2
M112 VDD ACTRCLK ACTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=10450 $Y=9420 $D=2
M113 DCTRCLKX 30 VDD VDD P12LL L=6E-08 W=5E-06 $X=10740 $Y=9420 $D=2
M114 VDD 30 DCTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=11030 $Y=9420 $D=2
M115 30 54 VDD VDD P12LL L=6E-08 W=3E-06 $X=11310 $Y=9420 $D=2
M116 58 22 VDD VDD P12LL L=6E-08 W=5E-06 $X=11900 $Y=9420 $D=2
M117 VDD 22 58 VDD P12LL L=6E-08 W=5E-06 $X=12190 $Y=9420 $D=2
M118 58 22 VDD VDD P12LL L=6E-08 W=5E-06 $X=12480 $Y=9420 $D=2
M119 VDD 22 58 VDD P12LL L=6E-08 W=5E-06 $X=12770 $Y=9420 $D=2
M120 56 58 VDD VDD P12LL L=6E-08 W=5E-06 $X=13640 $Y=9420 $D=2
M121 INTCLKX 57 56 VDD P12LL L=6E-08 W=5E-06 $X=13930 $Y=9420 $D=2
M122 56 57 INTCLKX VDD P12LL L=6E-08 W=5E-06 $X=14220 $Y=9420 $D=2
M123 VDD 58 56 VDD P12LL L=6E-08 W=5E-06 $X=14510 $Y=9420 $D=2
M124 56 58 VDD VDD P12LL L=6E-08 W=5E-06 $X=14800 $Y=9420 $D=2
M125 INTCLKX 57 56 VDD P12LL L=6E-08 W=5E-06 $X=15090 $Y=9420 $D=2
M126 56 57 INTCLKX VDD P12LL L=6E-08 W=5E-06 $X=15380 $Y=9420 $D=2
M127 VDD 58 56 VDD P12LL L=6E-08 W=5E-06 $X=15670 $Y=9420 $D=2
M128 57 59 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=15990 $Y=1440 $D=2
M129 VDD 59 57 VDD P12LL L=6E-08 W=1.4E-06 $X=16280 $Y=1440 $D=2
M130 59 58 VDD VDD P12LL L=6E-08 W=6E-07 $X=16570 $Y=2240 $D=2
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PX2                                                                 *
*******************************************************************************
.SUBCKT qspi_data_info_32_memPX2 VDD VSS PX[1] PX[0] A[0] CLK CLKX

M0 15 3 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=115 $Y=3520 $D=0
M1 PX[0] 4 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=115 $Y=10345 $D=0
M2 VSS 5 3 VSS N12LL L=6E-08 W=7E-07 $X=165 $Y=1550 $D=0
M3 8 CLKX 4 VSS N12LL L=6E-08 W=8.35E-07 $X=265 $Y=7855 $D=0
M4 VSS PX[0] 4 VSS N12LL L=6E-07 W=1.2E-07 $X=365 $Y=9535 $D=0
M5 8 VDD 15 VSS N12LL L=6E-08 W=7.5E-07 $X=405 $Y=3520 $D=0
M6 VSS 4 PX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=405 $Y=10345 $D=0
M7 5 6 VSS VSS N12LL L=6E-08 W=7E-07 $X=455 $Y=1550 $D=0
M8 4 CLKX 8 VSS N12LL L=6E-08 W=8.35E-07 $X=545 $Y=7855 $D=0
M9 16 VDD 8 VSS N12LL L=6E-08 W=7.5E-07 $X=695 $Y=3520 $D=0
M10 PX[0] 4 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=695 $Y=10345 $D=0
M11 8 CLKX 4 VSS N12LL L=6E-08 W=8.35E-07 $X=825 $Y=7855 $D=0
M12 VSS 3 16 VSS N12LL L=6E-08 W=7.5E-07 $X=985 $Y=3520 $D=0
M13 VSS 4 PX[0] VSS N12LL L=6E-08 W=7.5E-07 $X=985 $Y=10345 $D=0
M14 17 A[0] 6 VSS N12LL L=6E-08 W=4E-07 $X=1085 $Y=1550 $D=0
M15 18 5 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1275 $Y=3520 $D=0
M16 PX[1] 13 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1275 $Y=10345 $D=0
M17 VSS VDD 17 VSS N12LL L=3E-07 W=4E-07 $X=1325 $Y=1550 $D=0
M18 13 PX[1] VSS VSS N12LL L=6E-07 W=1.2E-07 $X=1355 $Y=9535 $D=0
M19 13 CLKX 14 VSS N12LL L=6E-08 W=8.35E-07 $X=1435 $Y=7855 $D=0
M20 14 VDD 18 VSS N12LL L=6E-08 W=7.5E-07 $X=1565 $Y=3520 $D=0
M21 VSS 13 PX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=1565 $Y=10345 $D=0
M22 14 CLKX 13 VSS N12LL L=6E-08 W=8.35E-07 $X=1715 $Y=7855 $D=0
M23 19 VDD 14 VSS N12LL L=6E-08 W=7.5E-07 $X=1855 $Y=3520 $D=0
M24 PX[1] 13 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=1855 $Y=10345 $D=0
M25 13 CLKX 14 VSS N12LL L=6E-08 W=8.35E-07 $X=1995 $Y=7855 $D=0
M26 VSS 5 19 VSS N12LL L=6E-08 W=7.5E-07 $X=2145 $Y=3520 $D=0
M27 VSS 13 PX[1] VSS N12LL L=6E-08 W=7.5E-07 $X=2145 $Y=10345 $D=0
M28 8 3 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=115 $Y=4770 $D=1
M29 PX[0] 4 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=115 $Y=11695 $D=1
M30 VDD 5 3 VDD P12LL L=6E-08 W=1.4E-06 $X=165 $Y=-450 $D=1
M31 8 CLK 4 VDD P12LL L=6E-08 W=8.3E-07 $X=265 $Y=6525 $D=1
M32 VDD VDD 8 VDD P12LL L=6E-08 W=7.5E-07 $X=405 $Y=4770 $D=1
M33 VDD 4 PX[0] VDD P12LL L=6E-08 W=1.75E-06 $X=405 $Y=11695 $D=1
M34 5 6 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=455 $Y=-450 $D=1
M35 4 CLK 8 VDD P12LL L=6E-08 W=8.3E-07 $X=545 $Y=6525 $D=1
M36 VDD PX[0] 4 VDD P12LL L=3E-07 W=1.2E-07 $X=615 $Y=14130 $D=1
M37 8 VDD VDD VDD P12LL L=6E-08 W=7.5E-07 $X=695 $Y=4770 $D=1
M38 PX[0] 4 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=695 $Y=11695 $D=1
M39 8 CLK 4 VDD P12LL L=6E-08 W=8.3E-07 $X=825 $Y=6525 $D=1
M40 VDD 3 8 VDD P12LL L=6E-08 W=7.5E-07 $X=985 $Y=4770 $D=1
M41 VDD 4 PX[0] VDD P12LL L=6E-08 W=1.75E-06 $X=985 $Y=11695 $D=1
M42 20 A[0] 6 VDD P12LL L=6E-08 W=4E-07 $X=1085 $Y=400 $D=1
M43 14 5 VDD VDD P12LL L=6E-08 W=7.5E-07 $X=1275 $Y=4770 $D=1
M44 PX[1] 13 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=1275 $Y=11695 $D=1
M45 13 PX[1] VDD VDD P12LL L=3E-07 W=1.2E-07 $X=1405 $Y=14130 $D=1
M46 VDD VSS 20 VDD P12LL L=1E-07 W=4E-07 $X=1425 $Y=400 $D=1
M47 13 CLK 14 VDD P12LL L=6E-08 W=8.3E-07 $X=1435 $Y=6525 $D=1
M48 VDD VDD 14 VDD P12LL L=6E-08 W=7.5E-07 $X=1565 $Y=4770 $D=1
M49 VDD 13 PX[1] VDD P12LL L=6E-08 W=1.75E-06 $X=1565 $Y=11695 $D=1
M50 14 CLK 13 VDD P12LL L=6E-08 W=8.3E-07 $X=1715 $Y=6525 $D=1
M51 14 VDD VDD VDD P12LL L=6E-08 W=7.5E-07 $X=1855 $Y=4770 $D=1
M52 PX[1] 13 VDD VDD P12LL L=6E-08 W=1.75E-06 $X=1855 $Y=11695 $D=1
M53 13 CLK 14 VDD P12LL L=6E-08 W=8.3E-07 $X=1995 $Y=6525 $D=1
M54 VDD 5 14 VDD P12LL L=6E-08 W=7.5E-07 $X=2145 $Y=4770 $D=1
M55 VDD 13 PX[1] VDD P12LL L=6E-08 W=1.75E-06 $X=2145 $Y=11695 $D=1
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TP_CLK                                                               *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTP_CLK VDD VSS ACTRCLK ACTRCLKX EMCLK INTCLKX SACK1 SACK4 CEN CLK FB

M0 VSS VSS VSS VSS N12LL L=1E-06 W=1E-06 $X=820 $Y=5625 $D=0
M1 VSS VSS VSS VSS N12LL L=1E-06 W=1E-06 $X=820 $Y=7600 $D=0
M2 VSS VSS VSS VSS N12LL L=1E-06 W=1E-06 $X=820 $Y=9340 $D=0
M3 35 CLK VSS VSS N12LL L=6E-08 W=4E-07 $X=1715 $Y=3545 $D=0
M4 79 35 VSS VSS N12LL L=6E-08 W=1E-06 $X=2365 $Y=3540 $D=0
M5 VSS VSS VSS VSS N12LL L=1E-06 W=1E-06 $X=2600 $Y=5625 $D=0
M6 VSS VSS VSS VSS N12LL L=1E-06 W=1E-06 $X=2600 $Y=7600 $D=0
M7 38 CEN 79 VSS N12LL L=6E-08 W=1E-06 $X=2605 $Y=3540 $D=0
M8 41 40 VSS VSS N12LL L=6E-08 W=1.25E-06 $X=2760 $Y=9475 $D=0
M9 VSS 40 41 VSS N12LL L=6E-08 W=1.25E-06 $X=3050 $Y=9475 $D=0
M10 VSS 51 38 VSS N12LL L=6E-07 W=1.2E-07 $X=3275 $Y=3830 $D=0
M11 40 FB VSS VSS N12LL L=6E-08 W=8E-07 $X=3340 $Y=9925 $D=0
M12 VSS 38 51 VSS N12LL L=6E-08 W=4E-07 $X=3920 $Y=3615 $D=0
M13 EMCLK 45 VSS VSS N12LL L=6E-08 W=6.05E-07 $X=4120 $Y=9995 $D=0
M14 44 51 VSS VSS N12LL L=6E-08 W=5E-07 $X=4210 $Y=3615 $D=0
M15 52 CLK 20 VSS N12LL L=6E-08 W=4E-06 $X=4280 $Y=4970 $D=0
M16 VSS 45 EMCLK VSS N12LL L=6E-08 W=6.05E-07 $X=4410 $Y=9995 $D=0
M17 VSS CLK 44 VSS N12LL L=6E-08 W=5E-07 $X=4500 $Y=3615 $D=0
M18 20 CLK 52 VSS N12LL L=6E-08 W=4E-06 $X=4570 $Y=4970 $D=0
M19 52 CLK 20 VSS N12LL L=6E-08 W=4E-06 $X=4860 $Y=4970 $D=0
M20 20 CLK 52 VSS N12LL L=6E-08 W=4E-06 $X=5150 $Y=4970 $D=0
M21 VSS 2 45 VSS N12LL L=2E-07 W=4E-07 $X=5165 $Y=10220 $D=0
M22 VSS 44 46 VSS N12LL L=6E-08 W=5E-07 $X=5190 $Y=3495 $D=0
M23 52 CLK 20 VSS N12LL L=6E-08 W=4E-06 $X=5440 $Y=4970 $D=0
M24 47 46 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=5540 $Y=3495 $D=0
M25 2 3 VSS VSS N12LL L=2E-07 W=4E-07 $X=5695 $Y=10220 $D=0
M26 VSS 46 47 VSS N12LL L=6E-08 W=7.5E-07 $X=5830 $Y=3495 $D=0
M27 52 47 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=6100 $Y=6125 $D=0
M28 VSS 47 52 VSS N12LL L=6E-08 W=2.5E-06 $X=6390 $Y=6125 $D=0
M29 VSS 50 3 VSS N12LL L=2E-07 W=4E-07 $X=6610 $Y=10220 $D=0
M30 52 47 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=6680 $Y=6125 $D=0
M31 VSS 47 52 VSS N12LL L=6E-08 W=2.5E-06 $X=6970 $Y=6125 $D=0
M32 VSS 53 21 VSS N12LL L=2E-07 W=4E-07 $X=7090 $Y=3435 $D=0
M33 50 20 VSS VSS N12LL L=6E-08 W=7E-07 $X=7100 $Y=9920 $D=0
M34 52 47 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=7260 $Y=6125 $D=0
M35 VSS 47 52 VSS N12LL L=6E-08 W=2.5E-06 $X=7550 $Y=6125 $D=0
M36 53 VSS VSS VSS N12LL L=2E-07 W=4E-07 $X=7580 $Y=3435 $D=0
M37 52 47 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=7840 $Y=6125 $D=0
M38 VSS 65 53 VSS N12LL L=2E-07 W=4E-07 $X=8070 $Y=3435 $D=0
M39 VSS 47 52 VSS N12LL L=6E-08 W=2.5E-06 $X=8130 $Y=6125 $D=0
M40 54 21 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=8420 $Y=6125 $D=0
M41 VSS 65 54 VSS N12LL L=6E-08 W=2.5E-06 $X=8710 $Y=6125 $D=0
M42 25 65 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=8975 $Y=3465 $D=0
M43 ACTRCLK 54 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=9000 $Y=6125 $D=0
M44 VSS 57 25 VSS N12LL L=6E-08 W=7.5E-07 $X=9265 $Y=3465 $D=0
M45 VSS 54 ACTRCLK VSS N12LL L=6E-08 W=2.5E-06 $X=9290 $Y=6125 $D=0
M46 25 57 VSS VSS N12LL L=6E-08 W=7.5E-07 $X=9555 $Y=3465 $D=0
M47 VSS 65 25 VSS N12LL L=6E-08 W=7.5E-07 $X=9845 $Y=3465 $D=0
M48 ACTRCLKX ACTRCLK VSS VSS N12LL L=6E-08 W=2.5E-06 $X=10160 $Y=6125 $D=0
M49 VSS ACTRCLK ACTRCLKX VSS N12LL L=6E-08 W=2.5E-06 $X=10450 $Y=6125 $D=0
M50 VSS 61 57 VSS N12LL L=2E-07 W=4E-07 $X=10555 $Y=3435 $D=0
M51 61 65 VSS VSS N12LL L=2E-07 W=4E-07 $X=11085 $Y=3435 $D=0
M52 SACK4 25 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=11320 $Y=6125 $D=0
M53 VSS 25 SACK4 VSS N12LL L=6E-08 W=2.5E-06 $X=11610 $Y=6125 $D=0
M54 65 20 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=11900 $Y=6125 $D=0
M55 VSS 65 20 VSS N12LL L=1E-06 W=1.2E-07 $X=11905 $Y=4325 $D=0
M56 VSS 20 65 VSS N12LL L=6E-08 W=2.5E-06 $X=12190 $Y=6125 $D=0
M57 65 20 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=12480 $Y=6125 $D=0
M58 VSS 20 65 VSS N12LL L=6E-08 W=2.5E-06 $X=12770 $Y=6125 $D=0
M59 SACK1 65 VSS VSS N12LL L=6E-08 W=2.5E-06 $X=13060 $Y=6125 $D=0
M60 VSS 65 SACK1 VSS N12LL L=6E-08 W=2.5E-06 $X=13350 $Y=6125 $D=0
M61 INTCLKX 65 VSS VSS N12LL L=6E-08 W=5E-06 $X=13640 $Y=3625 $D=0
M62 VSS 64 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=13930 $Y=3625 $D=0
M63 INTCLKX 64 VSS VSS N12LL L=6E-08 W=5E-06 $X=14220 $Y=3625 $D=0
M64 VSS 65 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=14510 $Y=3625 $D=0
M65 INTCLKX 65 VSS VSS N12LL L=6E-08 W=5E-06 $X=14800 $Y=3625 $D=0
M66 VSS 64 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=15090 $Y=3625 $D=0
M67 INTCLKX 64 VSS VSS N12LL L=6E-08 W=5E-06 $X=15380 $Y=3625 $D=0
M68 VSS 65 INTCLKX VSS N12LL L=6E-08 W=5E-06 $X=15670 $Y=3625 $D=0
M69 64 66 VSS VSS N12LL L=6E-08 W=7E-07 $X=15990 $Y=3625 $D=0
M70 VSS 66 64 VSS N12LL L=6E-08 W=7E-07 $X=16280 $Y=3625 $D=0
M71 66 65 VSS VSS N12LL L=6E-08 W=4E-07 $X=16570 $Y=3625 $D=0
M72 35 CLK VDD VDD P12LL L=6E-08 W=4E-07 $X=1715 $Y=2250 $D=2
M73 81 CLK VDD VDD P12LL L=6E-08 W=1E-06 $X=2365 $Y=1670 $D=2
M74 38 CEN 81 VDD P12LL L=6E-08 W=1E-06 $X=2605 $Y=1670 $D=2
M75 41 40 VDD VDD P12LL L=6E-08 W=1.24E-06 $X=2760 $Y=11385 $D=2
M76 VDD 51 38 VDD P12LL L=3E-07 W=1.2E-07 $X=2975 $Y=2435 $D=2
M77 VDD 40 41 VDD P12LL L=6E-08 W=1.24E-06 $X=3050 $Y=11385 $D=2
M78 40 FB VDD VDD P12LL L=6E-08 W=8E-07 $X=3340 $Y=11385 $D=2
M79 FB 50 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=3845 $Y=13320 $D=2
M80 VDD 38 51 VDD P12LL L=6E-08 W=8E-07 $X=3920 $Y=1870 $D=2
M81 EMCLK 45 VDD VDD P12LL L=6E-08 W=1.2E-06 $X=4120 $Y=11385 $D=2
M82 VDD 50 FB VDD P12LL L=6E-08 W=1.25E-06 $X=4135 $Y=13320 $D=2
M83 82 51 VDD VDD P12LL L=6E-08 W=1E-06 $X=4210 $Y=1670 $D=2
M84 VDD 45 EMCLK VDD P12LL L=6E-08 W=1.2E-06 $X=4410 $Y=11385 $D=2
M85 20 41 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=4425 $Y=13320 $D=2
M86 44 CLK 82 VDD P12LL L=6E-08 W=1E-06 $X=4500 $Y=1670 $D=2
M87 VDD 41 20 VDD P12LL L=6E-08 W=1.25E-06 $X=4715 $Y=13320 $D=2
M88 20 41 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5005 $Y=13320 $D=2
M89 VDD 2 45 VDD P12LL L=2E-07 W=6E-07 $X=5165 $Y=11385 $D=2
M90 VDD 44 46 VDD P12LL L=6E-08 W=1E-06 $X=5190 $Y=1800 $D=2
M91 VDD 41 20 VDD P12LL L=6E-08 W=1.25E-06 $X=5295 $Y=13320 $D=2
M92 47 46 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=5540 $Y=1300 $D=2
M93 20 41 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=5585 $Y=13320 $D=2
M94 2 3 VDD VDD P12LL L=2E-07 W=6E-07 $X=5695 $Y=11385 $D=2
M95 VDD 46 47 VDD P12LL L=6E-08 W=1.5E-06 $X=5830 $Y=1300 $D=2
M96 VDD 41 20 VDD P12LL L=6E-08 W=1.25E-06 $X=5875 $Y=13320 $D=2
M97 20 41 VDD VDD P12LL L=6E-08 W=1.25E-06 $X=6165 $Y=13320 $D=2
M98 VDD 41 20 VDD P12LL L=6E-08 W=1.25E-06 $X=6455 $Y=13320 $D=2
M99 VDD 50 3 VDD P12LL L=2E-07 W=6E-07 $X=6610 $Y=11385 $D=2
M100 VDD 53 21 VDD P12LL L=2E-07 W=4E-07 $X=7090 $Y=2165 $D=2
M101 50 20 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=7100 $Y=11385 $D=2
M102 83 VSS VDD VDD P12LL L=2E-07 W=8E-07 $X=7580 $Y=2165 $D=2
M103 53 65 83 VDD P12LL L=2E-07 W=8E-07 $X=8070 $Y=2165 $D=2
M104 84 21 54 VDD P12LL L=6E-08 W=5E-06 $X=8420 $Y=9420 $D=2
M105 VDD 65 84 VDD P12LL L=6E-08 W=5E-06 $X=8710 $Y=9420 $D=2
M106 55 65 VDD VDD P12LL L=6E-08 W=1.5E-06 $X=8975 $Y=1170 $D=2
M107 ACTRCLK 54 VDD VDD P12LL L=6E-08 W=5E-06 $X=9000 $Y=9420 $D=2
M108 25 57 55 VDD P12LL L=6E-08 W=1.5E-06 $X=9265 $Y=1170 $D=2
M109 VDD 54 ACTRCLK VDD P12LL L=6E-08 W=5E-06 $X=9290 $Y=9420 $D=2
M110 55 57 25 VDD P12LL L=6E-08 W=1.5E-06 $X=9555 $Y=1170 $D=2
M111 VDD 65 55 VDD P12LL L=6E-08 W=1.5E-06 $X=9845 $Y=1170 $D=2
M112 ACTRCLKX ACTRCLK VDD VDD P12LL L=6E-08 W=5E-06 $X=10160 $Y=9420 $D=2
M113 VDD ACTRCLK ACTRCLKX VDD P12LL L=6E-08 W=5E-06 $X=10450 $Y=9420 $D=2
M114 VDD 61 57 VDD P12LL L=2E-07 W=4E-07 $X=10555 $Y=2165 $D=2
M115 61 65 VDD VDD P12LL L=2E-07 W=4E-07 $X=11085 $Y=2165 $D=2
M116 SACK4 25 VDD VDD P12LL L=6E-08 W=5E-06 $X=11320 $Y=9420 $D=2
M117 VDD 25 SACK4 VDD P12LL L=6E-08 W=5E-06 $X=11610 $Y=9420 $D=2
M118 65 20 VDD VDD P12LL L=6E-08 W=5E-06 $X=11900 $Y=9420 $D=2
M119 20 65 VDD VDD P12LL L=2E-07 W=1.2E-07 $X=11945 $Y=2005 $D=2
M120 VDD 20 65 VDD P12LL L=6E-08 W=5E-06 $X=12190 $Y=9420 $D=2
M121 65 20 VDD VDD P12LL L=6E-08 W=5E-06 $X=12480 $Y=9420 $D=2
M122 VDD 20 65 VDD P12LL L=6E-08 W=5E-06 $X=12770 $Y=9420 $D=2
M123 SACK1 65 VDD VDD P12LL L=6E-08 W=5E-06 $X=13060 $Y=9420 $D=2
M124 VDD 65 SACK1 VDD P12LL L=6E-08 W=5E-06 $X=13350 $Y=9420 $D=2
M125 63 65 VDD VDD P12LL L=6E-08 W=5E-06 $X=13640 $Y=9420 $D=2
M126 INTCLKX 64 63 VDD P12LL L=6E-08 W=5E-06 $X=13930 $Y=9420 $D=2
M127 63 64 INTCLKX VDD P12LL L=6E-08 W=5E-06 $X=14220 $Y=9420 $D=2
M128 VDD 65 63 VDD P12LL L=6E-08 W=5E-06 $X=14510 $Y=9420 $D=2
M129 63 65 VDD VDD P12LL L=6E-08 W=5E-06 $X=14800 $Y=9420 $D=2
M130 INTCLKX 64 63 VDD P12LL L=6E-08 W=5E-06 $X=15090 $Y=9420 $D=2
M131 63 64 INTCLKX VDD P12LL L=6E-08 W=5E-06 $X=15380 $Y=9420 $D=2
M132 VDD 65 63 VDD P12LL L=6E-08 W=5E-06 $X=15670 $Y=9420 $D=2
M133 64 66 VDD VDD P12LL L=6E-08 W=1.4E-06 $X=15990 $Y=1440 $D=2
M134 VDD 66 64 VDD P12LL L=6E-08 W=1.4E-06 $X=16280 $Y=1440 $D=2
M135 66 65 VDD VDD P12LL L=6E-08 W=6E-07 $X=16570 $Y=2240 $D=2
.ENDS
***************************************
*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TPRWL_DEC                                                            *
*******************************************************************************
.SUBCKT qspi_data_info_32_memTPRWL_DEC VDD VSS RWL CLK CLKX RDE WLCKX

M0 23 VDD VSS VSS N12LL L=3E-07 W=4E-07 $X=485 $Y=285 $D=0
M1 7 5 VSS VSS N12LL L=6E-07 W=1.2E-07 $X=640 $Y=6180 $D=0
M2 VSS 5 3 VSS N12LL L=6E-08 W=4E-07 $X=665 $Y=4660 $D=0
M3 5 7 VSS VSS N12LL L=6E-08 W=4E-07 $X=965 $Y=4660 $D=0
M4 6 RDE 23 VSS N12LL L=6E-08 W=4E-07 $X=985 $Y=285 $D=0
M5 9 3 WLCKX VSS N12LL L=6E-08 W=5E-07 $X=1025 $Y=6960 $D=0
M6 RWL 9 VSS VSS N12LL L=6E-08 W=1E-06 $X=1025 $Y=10715 $D=0
M7 WLCKX 3 9 VSS N12LL L=6E-08 W=5E-07 $X=1315 $Y=6960 $D=0
M8 VSS 9 RWL VSS N12LL L=6E-08 W=1E-06 $X=1315 $Y=10715 $D=0
M9 9 3 WLCKX VSS N12LL L=6E-08 W=5E-07 $X=1605 $Y=6960 $D=0
M10 RWL 9 VSS VSS N12LL L=6E-08 W=1E-06 $X=1605 $Y=10715 $D=0
M11 VSS 6 12 VSS N12LL L=6E-08 W=4E-07 $X=1615 $Y=285 $D=0
M12 11 CLKX 7 VSS N12LL L=6E-08 W=1E-06 $X=1640 $Y=4800 $D=0
M13 WLCKX 3 9 VSS N12LL L=6E-08 W=5E-07 $X=1895 $Y=6960 $D=0
M14 VSS 9 RWL VSS N12LL L=6E-08 W=1E-06 $X=1895 $Y=10715 $D=0
M15 15 12 VSS VSS N12LL L=6E-08 W=4E-07 $X=1905 $Y=285 $D=0
M16 VSS 15 11 VSS N12LL L=6E-08 W=4E-07 $X=1940 $Y=4800 $D=0
M17 7 5 VDD VDD P12LL L=3E-07 W=1.2E-07 $X=540 $Y=2360 $D=1
M18 24 VSS VDD VDD P12LL L=1E-07 W=4E-07 $X=585 $Y=1520 $D=1
M19 VDD 5 3 VDD P12LL L=6E-08 W=8E-07 $X=665 $Y=3220 $D=1
M20 5 7 VDD VDD P12LL L=6E-08 W=8E-07 $X=965 $Y=3220 $D=1
M21 6 RDE 24 VDD P12LL L=6E-08 W=4E-07 $X=985 $Y=1520 $D=1
M22 9 5 WLCKX VDD P12LL L=6E-08 W=5E-07 $X=1025 $Y=8105 $D=1
M23 9 3 VDD VDD P12LL L=6E-08 W=5E-07 $X=1025 $Y=9075 $D=1
M24 RWL 9 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=1025 $Y=12445 $D=1
M25 WLCKX 5 9 VDD P12LL L=6E-08 W=5E-07 $X=1315 $Y=8105 $D=1
M26 VDD 3 9 VDD P12LL L=6E-08 W=5E-07 $X=1315 $Y=9075 $D=1
M27 VDD 9 RWL VDD P12LL L=6E-08 W=2.5E-06 $X=1315 $Y=12445 $D=1
M28 9 5 WLCKX VDD P12LL L=6E-08 W=5E-07 $X=1605 $Y=8105 $D=1
M29 9 3 VDD VDD P12LL L=6E-08 W=5E-07 $X=1605 $Y=9075 $D=1
M30 RWL 9 VDD VDD P12LL L=6E-08 W=2.5E-06 $X=1605 $Y=12445 $D=1
M31 VDD 6 12 VDD P12LL L=6E-08 W=8E-07 $X=1615 $Y=1465 $D=1
M32 11 CLK 7 VDD P12LL L=6E-08 W=1E-06 $X=1640 $Y=3020 $D=1
M33 WLCKX 5 9 VDD P12LL L=6E-08 W=5E-07 $X=1895 $Y=8105 $D=1
M34 VDD 3 9 VDD P12LL L=6E-08 W=5E-07 $X=1895 $Y=9075 $D=1
M35 VDD 9 RWL VDD P12LL L=6E-08 W=2.5E-06 $X=1895 $Y=12445 $D=1
M36 15 12 VDD VDD P12LL L=6E-08 W=8E-07 $X=1905 $Y=1465 $D=1
M37 VDD 15 11 VDD P12LL L=6E-08 W=8E-07 $X=1940 $Y=3220 $D=1
.ENDS
***************************************
*******************************************************************************
* MAIN CIRCUIT NETLIST:                                                       *
*                                                                             *
* BLOCK: qspi_data_info_32_mem                 *
                                                *
*******************************************************************************
.SUBCKT qspi_data_info_32_mem VDD VSS QA[31] QA[30]
+QA[29] QA[28] QA[27] QA[26] QA[25] QA[24] QA[23] QA[22] QA[21] QA[20]
+QA[19] QA[18] QA[17] QA[16] QA[15] QA[14] QA[13] QA[12] QA[11] QA[10]
+QA[9] QA[8] QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0]
+AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] 
+AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] 
+CENA CENB CLKA CLKB DB[31] 
+DB[30] DB[29] DB[28] DB[27] DB[26] DB[25] DB[24] DB[23] DB[22] DB[21] 
+DB[20] DB[19] DB[18] DB[17] DB[16] DB[15] DB[14] DB[13] DB[12] DB[11] 
+DB[10] DB[9] DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2] DB[1] 
+DB[0] 
XI4889 RDE VSS VDD qspi_data_info_32_mem_TIE_LOW_X2
XI4888_0 TIE_LOW VSS VDD qspi_data_info_32_mem_TIE_LOW_X1
XI4888_1 TIE_HIGH VSS VDD qspi_data_info_32_mem_TIE_HIGH_X1
XI15 VDD VSS FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0]
+AB[0] AB[1] AB[2] ACTRCLKB ACTRCLKXB INTCLKXB qspi_data_info_32_memFPREDEC
XI9 VDD VSS FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0]
+AA[0] AA[1] AA[2] ACTRCLKA ACTRCLKXA INTCLKXA qspi_data_info_32_memFPREDEC
XI6 VDD VSS PXAA[3] PXAA[2] PXAA[1] PXAA[0] AA[3] AA[4] ACTRCLKA ACTRCLKXA RDE  qspi_data_info_32_memPXA
XI1 VDD VSS PXAB[3] PXAB[2] PXAB[1] PXAB[0] AB[3] AB[4] ACTRCLKB ACTRCLKXB RDE  qspi_data_info_32_memPXA
XI8 VDD VSS PXBA[1] PXBA[0] AA[5] ACTRCLKA ACTRCLKXA qspi_data_info_32_memPX2
XI14 VDD VSS PXBB[1] PXBB[0] AB[5] ACTRCLKB ACTRCLKXB qspi_data_info_32_memPX2
XI21 VDD VSS DBLA EMCLKA SOPA[5] SOPA[4] SOPA[3] SOPA[2] SOPA[1] SOPA[0]
+qspi_data_info_32_memTP_DISCHARGECELLS
XI19 VDD VSS QA[15] QA[14] QA[13] QA[12] QA[11] QA[10] QA[9] QA[8] 
+QA[7] QA[6] QA[5] QA[4] QA[3] QA[2] QA[1] QA[0] 
+BWENB[15] BWENB[14] BWENB[13] BWENB[12] BWENB[11] BWENB[10] BWENB[9] BWENB[8] 
+BWENB[7] BWENB[6] BWENB[5] BWENB[4] BWENB[3] BWENB[2] BWENB[1] BWENB[0] 
+SACK1 SACK4 DCTRCLKW DCTRCLKXW
+DB[15] DB[14] DB[13] DB[12] DB[11] DB[10] DB[9] 
+DB[8] DB[7] DB[6] DB[5] DB[4] DB[3] DB[2] DB[1] 
+DB[0] INTCLKXB VSS RWLA[1] VSS RWLB[1] WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+qspi_data_info_32_memTPRF_X64Y1D16
XI18 VDD VSS QA[31] QA[30] QA[29] QA[28] QA[27] QA[26] QA[25] QA[24] 
+QA[23] QA[22] QA[21] QA[20] QA[19] QA[18] QA[17] QA[16] 
+BWENB[31] BWENB[30] BWENB[29] BWENB[28] BWENB[27] BWENB[26] BWENB[25] BWENB[24] 
+BWENB[23] BWENB[22] BWENB[21] BWENB[20] BWENB[19] BWENB[18] BWENB[17] BWENB[16] 
+SACK1 SACK4 DCTRCLKW DCTRCLKXW DBLA DB[31] 
+DB[30] DB[29] DB[28] DB[27] DB[26] DB[25] DB[24] DB[23] DB[22] DB[21] 
+DB[20] DB[19] DB[18] DB[17] DB[16] INTCLKXB VSS RWLA[1] VSS RWLB[1] WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+qspi_data_info_32_memTPRF_X64Y1D16_ST
XI23 VDD VSS AA[5] AA[4] AA[3] AA[2] AA[1] AA[0] 
+CENA CLKA qspi_data_info_32_memESDA5W
XI12 VDD VSS AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] 
+CENB CLKB RDE  qspi_data_info_32_memESDA5R
XI22 VDD VSS SOPA[5] SOPA[4] SOPA[3] SOPA[2] SOPA[1] SOPA[0] TIE_LOW TIE_HIGH TIE_HIGH qspi_data_info_32_memOPDEC
XI16 VDD VSS WLB[63] WLB[62] WLB[61] WLB[60]
+WLB[59] WLB[58] WLB[57] WLB[56] WLB[55] WLB[54] WLB[53] WLB[52] WLB[51] WLB[50]
+WLB[49] WLB[48] WLB[47] WLB[46] WLB[45] WLB[44] WLB[43] WLB[42] WLB[41] WLB[40]
+WLB[39] WLB[38] WLB[37] WLB[36] WLB[35] WLB[34] WLB[33] WLB[32] WLB[31] WLB[30]
+WLB[29] WLB[28] WLB[27] WLB[26] WLB[25] WLB[24] WLB[23] WLB[22] WLB[21] WLB[20]
+WLB[19] WLB[18] WLB[17] WLB[16] WLB[15] WLB[14] WLB[13] WLB[12] WLB[11] WLB[10]
+WLB[9] WLB[8] WLB[7] WLB[6] WLB[5] WLB[4] WLB[3] WLB[2] WLB[1] WLB[0]
+FCKXB[7] FCKXB[6] FCKXB[5] FCKXB[4] FCKXB[3] FCKXB[2] FCKXB[1] FCKXB[0]
+PXAB[3] PXAB[2] PXAB[1] PXAB[0] PXBB[1] PXBB[0] VDD qspi_data_info_32_memXDEC8
XI17 VDD VSS WLA[63] WLA[62] WLA[61] WLA[60]
+WLA[59] WLA[58] WLA[57] WLA[56] WLA[55] WLA[54] WLA[53] WLA[52] WLA[51] WLA[50]
+WLA[49] WLA[48] WLA[47] WLA[46] WLA[45] WLA[44] WLA[43] WLA[42] WLA[41] WLA[40]
+WLA[39] WLA[38] WLA[37] WLA[36] WLA[35] WLA[34] WLA[33] WLA[32] WLA[31] WLA[30]
+WLA[29] WLA[28] WLA[27] WLA[26] WLA[25] WLA[24] WLA[23] WLA[22] WLA[21] WLA[20]
+WLA[19] WLA[18] WLA[17] WLA[16] WLA[15] WLA[14] WLA[13] WLA[12] WLA[11] WLA[10]
+WLA[9] WLA[8] WLA[7] WLA[6] WLA[5] WLA[4] WLA[3] WLA[2] WLA[1] WLA[0]
+FCKXA[7] FCKXA[6] FCKXA[5] FCKXA[4] FCKXA[3] FCKXA[2] FCKXA[1] FCKXA[0]
+PXAA[3] PXAA[2] PXAA[1] PXAA[0] PXBA[1] PXBA[0] VDD qspi_data_info_32_memXDEC8
XI10 VDD VSS ACTRCLKB ACTRCLKXB DCTRCLKW DCTRCLKXW INTCLKXB CENB CLKB qspi_data_info_32_memTP_CLKW
XI5 VDD VSS ACTRCLKA ACTRCLKXA EMCLKA INTCLKXA SACK1 SACK4 CENA CLKA DBLA qspi_data_info_32_memTP_CLK
XI4 VDD VSS RWLA[1] ACTRCLKA ACTRCLKXA RDE INTCLKXA qspi_data_info_32_memTPRWL_DEC
XI11 VDD VSS RWLB[1] ACTRCLKB ACTRCLKXB RDE INTCLKXB qspi_data_info_32_memTPRWL_DEC
.ENDS qspi_data_info_32_mem
